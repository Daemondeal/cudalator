module file1;
    int x;

    always_comb x = 2;
endmodule

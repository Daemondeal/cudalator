module file2;
    file1 file1_1_i();
    file1 file1_2_i();
endmodule

module int_adder (
    input int a,
    input int b,
    output int sum
);
assign sum = a + b;

endmodule : int_adder

module simple (
    output logic [7:0] value
);

endmodule : simple

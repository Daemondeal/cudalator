module first(input x, output z);
logic x;
logic z;

assign z = ~x;

endmodule

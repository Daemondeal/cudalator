module second;

logic x;
logic z;

first first_i (x, z);

endmodule

//# 35 inputs
//# 49 outputs
//# 179 D-type flipflops
//# 1775 inverters
//# 1004 gates (0 ANDs + 0 NANDs + 239 ORs + 765 NORs)

module dff (CK,Q,D);
input CK,D;
output Q;
reg Q;
always @ (posedge CK)
  Q <= D;
endmodule

module s5378(CK,n3065gat,n3066gat,n3067gat,n3068gat,n3069gat,n3070gat,
  n3071gat,
  n3072gat,n3073gat,n3074gat,n3075gat,n3076gat,n3077gat,n3078gat,n3079gat,
  n3080gat,n3081gat,n3082gat,n3083gat,n3084gat,n3085gat,n3086gat,n3087gat,
  n3088gat,n3089gat,n3090gat,n3091gat,n3092gat,n3093gat,n3094gat,n3095gat,
  n3097gat,n3098gat,n3099gat,n3100gat,n3104gat,n3105gat,n3106gat,n3107gat,
  n3108gat,n3109gat,n3110gat,n3111gat,n3112gat,n3113gat,n3114gat,n3115gat,
  n3116gat,n3117gat,n3118gat,n3119gat,n3120gat,n3121gat,n3122gat,n3123gat,
  n3124gat,n3125gat,n3126gat,n3127gat,n3128gat,n3129gat,n3130gat,n3131gat,
  n3132gat,n3133gat,n3134gat,n3135gat,n3136gat,n3137gat,n3138gat,n3139gat,
  n3140gat,n3141gat,n3142gat,n3143gat,n3144gat,n3145gat,n3146gat,n3147gat,
  n3148gat,n3149gat,n3150gat,n3151gat,n3152gat);
input CK,n3065gat,n3066gat,n3067gat,n3068gat,n3069gat,n3070gat,
  n3071gat,n3072gat,
  n3073gat,n3074gat,n3075gat,n3076gat,n3077gat,n3078gat,n3079gat,n3080gat,
  n3081gat,n3082gat,n3083gat,n3084gat,n3085gat,n3086gat,n3087gat,n3088gat,
  n3089gat,n3090gat,n3091gat,n3092gat,n3093gat,n3094gat,n3095gat,n3097gat,
  n3098gat,n3099gat,n3100gat;
output n3104gat,n3105gat,n3106gat,n3107gat,n3108gat,n3109gat,n3110gat,n3111gat,
  n3112gat,n3113gat,n3114gat,n3115gat,n3116gat,n3117gat,n3118gat,n3119gat,
  n3120gat,n3121gat,n3122gat,n3123gat,n3124gat,n3125gat,n3126gat,n3127gat,
  n3128gat,n3129gat,n3130gat,n3131gat,n3132gat,n3133gat,n3134gat,n3135gat,
  n3136gat,n3137gat,n3138gat,n3139gat,n3140gat,n3141gat,n3142gat,n3143gat,
  n3144gat,n3145gat,n3146gat,n3147gat,n3148gat,n3149gat,n3150gat,n3151gat,
  n3152gat;

  wire n673gat,n2897gat,n398gat,n2782gat,n402gat,n2790gat,n919gat,n2670gat,
    n846gat,n2793gat,n394gat,n703gat,n722gat,n726gat,n2510gat,n748gat,n271gat,
    n2732gat,n160gat,n2776gat,n337gat,n2735gat,n842gat,n2673gat,n341gat,
    n2779gat,n2522gat,n43gat,n2472gat,n1620gat,n2319gat,n2470gat,n1821gat,
    n1827gat,n1825gat,n2029gat,n1816gat,n1829gat,n2027gat,n283gat,n165gat,
    n279gat,n1026gat,n275gat,n2476gat,n55gat,n1068gat,n2914gat,n957gat,
    n2928gat,n861gat,n2927gat,n1294gat,n2896gat,n1241gat,n2922gat,n1298gat,
    n865gat,n2894gat,n1080gat,n2921gat,n1148gat,n2895gat,n2468gat,n933gat,
    n618gat,n491gat,n622gat,n626gat,n834gat,n3064gat,n707gat,n3055gat,n838gat,
    n3063gat,n830gat,n3062gat,n614gat,n3056gat,n2526gat,n504gat,n680gat,
    n2913gat,n816gat,n2920gat,n580gat,n2905gat,n824gat,n3057gat,n820gat,
    n3059gat,n883gat,n3058gat,n584gat,n2898gat,n684gat,n3060gat,n699gat,
    n3061gat,n2464gat,n567gat,n2399gat,n3048gat,n2343gat,n3049gat,n2203gat,
    n3051gat,n2562gat,n3047gat,n2207gat,n3050gat,n2626gat,n3040gat,n2490gat,
    n3044gat,n2622gat,n3042gat,n2630gat,n3037gat,n2543gat,n3041gat,n2102gat,
    n1606gat,n1880gat,n3052gat,n1763gat,n1610gat,n2155gat,n1858gat,n1035gat,
    n2918gat,n1121gat,n2952gat,n1072gat,n2919gat,n1282gat,n2910gat,n1226gat,
    n2907gat,n931gat,n2911gat,n1135gat,n2912gat,n1045gat,n2909gat,n1197gat,
    n2908gat,n2518gat,n2971gat,n667gat,n2904gat,n659gat,n2891gat,n553gat,
    n2903gat,n777gat,n2915gat,n561gat,n2901gat,n366gat,n2890gat,n322gat,
    n2888gat,n318gat,n2887gat,n314gat,n2886gat,n2599gat,n3010gat,n2588gat,
    n3016gat,n2640gat,n3054gat,n2658gat,n2579gat,n2495gat,n3036gat,n2390gat,
    n3034gat,n2270gat,n3031gat,n2339gat,n3035gat,n2502gat,n2646gat,n2634gat,
    n3053gat,n2506gat,n2613gat,n1834gat,n1625gat,n1767gat,n1626gat,n2084gat,
    n1603gat,n2143gat,n2541gat,n2061gat,n2557gat,n2139gat,n2487gat,n1899gat,
    n2532gat,n1850gat,n2628gat,n2403gat,n2397gat,n2394gat,n2341gat,n2440gat,
    n2560gat,n2407gat,n2205gat,n2347gat,n2201gat,n1389gat,n1793gat,n2021gat,
    n1781gat,n1394gat,n1516gat,n1496gat,n1392gat,n2091gat,n1685gat,n1332gat,
    n1565gat,n1740gat,n1330gat,n2179gat,n1945gat,n2190gat,n2268gat,n2135gat,
    n2337gat,n2262gat,n2388gat,n2182gat,n1836gat,n1433gat,n2983gat,n1316gat,
    n1431gat,n1363gat,n1314gat,n1312gat,n1361gat,n1775gat,n1696gat,n1871gat,
    n2009gat,n2592gat,n1773gat,n1508gat,n1636gat,n1678gat,n1712gat,n2309gat,
    n3000gat,n2450gat,n2307gat,n2446gat,n2661gat,n2095gat,n827gat,n2176gat,
    n2093gat,n2169gat,n2174gat,n2454gat,n2163gat,n2040gat,n1777gat,n2044gat,
    n2015gat,n2037gat,n2042gat,n2025gat,n2017gat,n2099gat,n2023gat,n2266gat,
    n2493gat,n2033gat,n2035gat,n2110gat,n2031gat,n2125gat,n2108gat,n2121gat,
    n2123gat,n2117gat,n2119gat,n1975gat,n2632gat,n2644gat,n2638gat,n156gat,
    n612gat,n152gat,n705gat,n331gat,n822gat,n388gat,n881gat,n463gat,n818gat,
    n327gat,n682gat,n384gat,n697gat,n256gat,n836gat,n470gat,n828gat,n148gat,
    n832gat,n2458gat,n2590gat,n2514gat,n2456gat,n1771gat,n1613gat,n1336gat,
    n1391gat,n1748gat,n1927gat,n1675gat,n1713gat,n1807gat,n1717gat,n1340gat,
    n1567gat,n1456gat,n1564gat,n1525gat,n1632gat,n1462gat,n1915gat,n1596gat,
    n1800gat,n1588gat,n1593gat,II1,n2717gat,n2715gat,II5,n2725gat,n2723gat,
    n296gat,n421gat,II11,n2768gat,II14,n2767gat,n373gat,II18,n2671gat,n2669gat,
    II23,n2845gat,n2844gat,II27,n2668gat,II30,n2667gat,n856gat,II44,n672gat,
    II47,n2783gat,II50,n396gat,II62,n2791gat,II65,II76,n401gat,n1645gat,
    n1499gat,II81,II92,n918gat,n1553gat,n1616gat,II97,n2794gat,II100,II111,
    n845gat,n1559gat,n1614gat,n1643gat,n1641gat,n1651gat,n1642gat,n1562gat,
    n1556gat,n1560gat,n1557gat,n1640gat,n1639gat,n1566gat,n1605gat,n1554gat,
    n1555gat,n1722gat,n1558gat,n392gat,II149,n702gat,n1319gat,n1256gat,n720gat,
    II171,n725gat,n1447gat,n1117gat,n1627gat,n1618gat,II178,n721gat,n1380gat,
    n1114gat,n1628gat,n1621gat,n701gat,n1446gat,n1318gat,n1705gat,n1619gat,
    n1706gat,n1622gat,II192,n2856gat,n2854gat,II196,n1218gat,II199,n2861gat,
    n2859gat,II203,n1219gat,II206,n2864gat,n2862gat,II210,n1220gat,II214,
    n2860gat,II217,n1221gat,II220,n2863gat,II223,n1222gat,II227,n2855gat,II230,
    n1223gat,n640gat,n1213gat,II237,n753gat,II240,n2716gat,II243,n2869gat,
    n2867gat,II248,n2868gat,II253,n2906gat,n754gat,II256,n2724gat,II259,
    n2728gat,n2726gat,II264,n2727gat,n422gat,n2889gat,II270,n755gat,n747gat,
    II275,n756gat,II278,n757gat,II282,n758gat,n2508gat,II297,n2733gat,II300,
    II311,n270gat,II314,n263gat,II317,n2777gat,II320,II331,n159gat,II334,
    n264gat,II337,n2736gat,II340,II351,n336gat,II354,n265gat,n158gat,II359,
    n266gat,n335gat,II363,n267gat,n269gat,II368,n268gat,n41gat,n258gat,II375,
    n48gat,II378,n1018gat,II381,n2674gat,II384,II395,n841gat,II398,n1019gat,
    II401,n1020gat,n840gat,II406,n1021gat,II409,n1022gat,n724gat,II414,
    n1023gat,II420,n1013gat,n49gat,II423,n2780gat,II426,II437,n340gat,II440,
    n480gat,II443,n481gat,II446,n393gat,II449,n482gat,II453,n483gat,II456,
    n484gat,n339gat,II461,n485gat,n42gat,n475gat,II468,n50gat,n162gat,II473,
    n51gat,II476,n52gat,II480,n53gat,n2520gat,n1448gat,n1376gat,n1701gat,
    n1617gat,n1379gat,n1377gat,n1615gat,n1624gat,n1500gat,n1113gat,n1503gat,
    n1501gat,n1779gat,n1623gat,II509,n2730gat,II512,n2729gat,n2317gat,n1819gat,
    n1823gat,n1817gat,II572,n1828gat,II576,n2851gat,II579,n2850gat,II583,
    n2786gat,n2785gat,n92gat,n637gat,n529gat,n293gat,n361gat,II591,n2722gat,
    II594,n2721gat,n297gat,II606,n282gat,II609,n172gat,II620,n164gat,II623,
    n173gat,II634,n278gat,II637,n174gat,n163gat,II642,n175gat,n277gat,II646,
    n176gat,n281gat,II651,n177gat,n54gat,n167gat,II658,n60gat,II661,n911gat,
    II672,n1025gat,II675,n912gat,II678,n913gat,n1024gat,II683,n914gat,n917gat,
    II687,n915gat,n844gat,II692,n916gat,II698,n906gat,n61gat,II709,n274gat,
    II712,n348gat,II715,n349gat,II718,n397gat,II721,n350gat,n400gat,II726,
    n351gat,II729,n352gat,n273gat,II734,n353gat,n178gat,n343gat,II741,n62gat,
    n66gat,II746,n63gat,II749,n64gat,II753,n65gat,n2474gat,II768,n2832gat,
    II771,n2831gat,n2731gat,II776,n2719gat,n2718gat,II790,n1067gat,II793,
    n949gat,II796,n2839gat,n2838gat,n2775gat,II812,n956gat,II815,n950gat,II818,
    n2712gat,n2711gat,n2734gat,II834,n860gat,II837,n951gat,n955gat,II842,
    n952gat,n859gat,II846,n953gat,n1066gat,II851,n954gat,n857gat,n944gat,II858,
    n938gat,n2792gat,II863,n2847gat,n2846gat,II877,n1293gat,II880,n1233gat,
    n2672gat,II885,n2853gat,n2852gat,II899,n1240gat,II902,n1234gat,II913,
    n1297gat,II916,n1235gat,n1239gat,II921,n1236gat,n1296gat,II925,n1237gat,
    n1292gat,II930,n1238gat,II936,n1228gat,n939gat,n2778gat,II941,n2837gat,
    n2836gat,II955,n864gat,II958,n1055gat,n2789gat,II963,n2841gat,n2840gat,
    II977,n1079gat,II980,n1056gat,n2781gat,II985,n2843gat,n2842gat,II999,
    n1147gat,II1002,n1057gat,n1078gat,II1007,n1058gat,n1146gat,II1011,n1059gat,
    n863gat,II1016,n1060gat,n928gat,n1050gat,II1023,n940gat,n858gat,II1028,
    n941gat,II1031,n942gat,II1035,n943gat,n2466gat,n2720gat,n740gat,n2784gat,
    n743gat,n746gat,n294gat,n360gat,n374gat,n616gat,II1067,n501gat,n489gat,
    II1079,n502gat,II1082,n617gat,II1085,n499gat,II1088,n490gat,II1091,n500gat,
    n620gat,II1103,n738gat,n624gat,II1115,n737gat,II1118,n621gat,II1121,
    n733gat,II1124,n625gat,II1127,n735gat,II1138,n833gat,II1141,n714gat,II1152,
    n706gat,II1155,n715gat,II1166,n837gat,II1169,n716gat,II1174,n717gat,II1178,
    n718gat,II1183,n719gat,n515gat,n709gat,II1190,n509gat,II1201,n829gat,
    II1204,n734gat,II1209,n736gat,II1216,n728gat,n510gat,II1227,n613gat,II1230,
    n498gat,II1236,n503gat,n404gat,n493gat,II1243,n511gat,n405gat,II1248,
    n512gat,II1251,n513gat,II1255,n514gat,n2524gat,n17gat,n564gat,n79gat,
    n86gat,n219gat,n78gat,n563gat,II1278,n289gat,n179gat,n287gat,n188gat,
    n288gat,n72gat,n181gat,n111gat,n182gat,II1302,n679gat,II1305,n808gat,
    II1319,n815gat,II1322,n809gat,II1336,n579gat,II1339,n810gat,n814gat,II1344,
    n811gat,n578gat,II1348,n812gat,n678gat,II1353,n813gat,n677gat,n803gat,
    II1360,n572gat,II1371,n823gat,II1374,n591gat,II1385,n819gat,II1388,n592gat,
    II1399,n882gat,II1402,n593gat,II1407,n594gat,II1411,n595gat,II1416,n596gat,
    II1422,n586gat,n573gat,II1436,n583gat,II1439,n691gat,II1450,n683gat,II1453,
    n692gat,II1464,n698gat,II1467,n693gat,II1472,n694gat,II1476,n695gat,
    n582gat,II1481,n696gat,n456gat,n686gat,II1488,n574gat,n565gat,II1493,
    n575gat,II1496,n576gat,II1500,n577gat,n2462gat,n2665gat,II1516,n2596gat,
    n189gat,n286gat,n194gat,n187gat,n21gat,n15gat,II1538,n2398gat,n2353gat,
    II1550,n2342gat,n2284gat,n2354gat,n2356gat,n2214gat,n2286gat,II1585,
    n2624gat,II1606,n2489gat,II1617,n2621gat,n2533gat,n2534gat,II1630,n2629gat,
    n2486gat,n2429gat,n2432gat,n2430gat,II1655,n2101gat,n1693gat,II1667,
    n1879gat,n1698gat,n1934gat,n1543gat,II1683,n1762gat,n1673gat,n2989gat,
    II1698,n2154gat,n2488gat,II1703,n2625gat,n2530gat,n2531gat,II1708,n2542gat,
    n2482gat,n2426gat,n2480gat,n2153gat,n2355gat,II1719,n2561gat,n2443gat,
    n2289gat,II1724,n2148gat,II1734,n855gat,n759gat,II1749,n1034gat,II1752,
    n1189gat,n1075gat,II1766,n1120gat,II1769,n1190gat,n760gat,II1783,n1071gat,
    II1786,n1191gat,n1119gat,II1791,n1192gat,n1070gat,II1795,n1193gat,n1033gat,
    II1800,n1194gat,n1183gat,n1184gat,II1807,n1274gat,n644gat,n1280gat,n641gat,
    II1833,n1225gat,II1837,n1281gat,n1224gat,II1843,n2970gat,n1275gat,n761gat,
    II1857,n930gat,II1860,n1206gat,n762gat,II1874,n1134gat,II1877,n1207gat,
    n643gat,II1891,n1044gat,II1894,n1208gat,n1133gat,II1899,n1209gat,n1043gat,
    II1903,n1210gat,n929gat,II1908,n1211gat,n1268gat,n1201gat,II1915,n1276gat,
    n1329gat,II1920,n1277gat,II1923,n1278gat,II1927,n1279gat,n1284gat,n1269gat,
    n642gat,n1195gat,II1947,n1196gat,n2516gat,II1961,n3017gat,n851gat,n853gat,
    n1725gat,n664gat,n852gat,n854gat,II1981,n666gat,n368gat,II1996,n658gat,
    II1999,n784gat,n662gat,II2014,n552gat,II2017,n785gat,n661gat,II2032,
    n776gat,II2035,n786gat,n551gat,II2040,n787gat,n775gat,II2044,n788gat,
    n657gat,II2049,n789gat,n35gat,n779gat,II2056,n125gat,n558gat,n559gat,
    n371gat,II2084,n365gat,II2088,n560gat,n364gat,II2094,n2876gat,n126gat,
    n663gat,II2109,n321gat,II2112,n226gat,n370gat,II2127,n317gat,II2130,
    n227gat,n369gat,II2145,n313gat,II2148,n228gat,n316gat,II2153,n229gat,
    n312gat,II2157,n230gat,n320gat,II2162,n231gat,n34gat,n221gat,II2169,
    n127gat,n133gat,II2174,n128gat,II2177,n129gat,II2181,n130gat,n665gat,
    n1601gat,n120gat,n2597gat,n2595gat,n2594gat,n2586gat,II2213,n2573gat,
    II2225,n2574gat,II2228,n2575gat,II2232,n2639gat,II2235,n2576gat,II2238,
    n2577gat,II2242,n2578gat,II2248,n2568gat,n2582gat,II2251,n2206gat,II2254,
    n2414gat,II2257,n2415gat,II2260,n2202gat,II2263,n2416gat,II2268,n2417gat,
    II2271,n2418gat,II2275,n2419gat,II2281,n2409gat,n2585gat,n2656gat,II2316,
    n2389gat,II2319,n2494gat,II2324,n3014gat,n2649gat,II2344,n2338gat,II2349,
    n2269gat,II2354,n2880gat,n2652gat,n2500gat,n2620gat,n2612gat,II2372,
    n2606gat,II2376,n2607gat,n2540gat,II2380,n2608gat,n2536gat,II2385,n2609gat,
    II2389,n2610gat,II2394,n2611gat,II2400,n2601gat,n2616gat,II2403,n2550gat,
    II2414,n2633gat,II2417,n2551gat,II2420,n2552gat,II2425,n2553gat,II2428,
    n2554gat,II2433,n2555gat,II2439,n2545gat,n2619gat,n2504gat,n2660gat,
    n2655gat,n1528gat,n2293gat,n1523gat,n2219gat,n1592gat,n1529gat,n2666gat,
    n1704gat,n2422gat,n3013gat,n2290gat,n2081gat,n2218gat,n2285gat,n2359gat,
    n2358gat,n1414gat,n1415gat,n566gat,n1480gat,n2292gat,n1301gat,n1416gat,
    n1150gat,n873gat,n2011gat,n2306gat,n1478gat,n1481gat,n875gat,n1410gat,
    n2357gat,n876gat,n1347gat,n1160gat,n1484gat,n1084gat,n983gat,n1482gat,
    n2363gat,n1157gat,n1483gat,n985gat,n1530gat,n2364gat,n1307gat,n1308gat,
    n1085gat,n1479gat,n2291gat,n1348gat,n1349gat,n2217gat,n1591gat,n2223gat,
    n1437gat,n1438gat,n1832gat,n1765gat,n1878gat,n1442gat,n1831gat,n1444gat,
    n1378gat,n2975gat,n1322gat,n2974gat,n1439gat,n1486gat,n1370gat,n1426gat,
    n1369gat,n2966gat,n1366gat,n1365gat,n1374gat,n2979gat,n2162gat,n2220gat,
    n1450gat,n1423gat,n1427gat,n1608gat,n2082gat,n1449gat,n1494gat,n1590gat,
    n1248gat,n2954gat,n1418gat,n1417gat,n1306gat,n2964gat,n1353gat,n1419gat,
    n1247gat,n2958gat,n1355gat,n1422gat,n1300gat,n2963gat,n1487gat,n1485gat,
    n1164gat,n2953gat,n1356gat,n1354gat,n1436gat,n1435gat,n1106gat,n2949gat,
    n1425gat,n1421gat,n1105gat,n2934gat,n1424gat,n1420gat,n1309gat,n2959gat,
    II2672,n2142gat,n1788gat,II2684,n2060gat,n1786gat,II2696,n2138gat,n1839gat,
    n1897gat,n1884gat,n1848gat,n1783gat,n1548gat,II2721,n1719gat,n2137gat,
    n1633gat,n2059gat,n1785gat,II2731,n1849gat,n1784gat,n1716gat,II2736,
    n1635gat,n2401gat,n1989gat,n2392gat,n1918gat,II2771,n2439gat,n1986gat,
    n1866gat,n1865gat,II2785,n2406gat,n2216gat,n2345gat,n1988gat,n1735gat,
    n1861gat,n1387gat,n1694gat,II2813,n1780gat,n2019gat,n1549gat,II2832,
    n1551gat,II2837,n2346gat,n2152gat,n2405gat,n2351gat,II2843,n2402gat,
    n2212gat,II2847,n2393gat,n1991gat,n1665gat,n1666gat,n1517gat,n1578gat,
    II2873,n1495gat,n1604gat,II2885,n2090gat,n1550gat,II2890,n1552gat,n1738gat,
    II2915,n1739gat,n1925gat,n1920gat,n1917gat,n1921gat,n2141gat,n1787gat,
    II2926,n1859gat,n1922gat,n1798gat,II2935,n1743gat,n1923gat,n1864gat,
    n1690gat,II2953,n2178gat,n1661gat,n1660gat,n1572gat,n1576gat,n2438gat,
    n2283gat,n1520gat,n1582gat,n1580gat,n1577gat,n1990gat,n2988gat,II2978,
    n2189gat,II2989,n2134gat,II3000,n2261gat,n2128gat,n2129gat,n1695gat,II3016,
    n2181gat,II3056,n1311gat,n1707gat,n1659gat,n2987gat,n1515gat,n1521gat,
    n1736gat,n1737gat,n1658gat,n1724gat,n1732gat,n1662gat,n1663gat,n1656gat,
    n1655gat,n1670gat,n1667gat,n1569gat,n1570gat,n1568gat,n1575gat,n1727gat,
    n1728gat,n1797gat,n1801gat,n1730gat,n1731gat,n1561gat,n1571gat,n1668gat,
    n1734gat,n1742gat,n1671gat,n1669gat,n1652gat,n1657gat,n1648gat,n1729gat,
    n1790gat,n1726gat,n2004gat,n1929gat,n1869gat,II3143,n2591gat,n1584gat,
    n1714gat,II3149,n1718gat,II3163,n1507gat,n1396gat,n1401gat,II3168,n1393gat,
    n1409gat,n1476gat,II3174,n1898gat,n1838gat,II3179,II3191,n1677gat,n2000gat,
    n1412gat,n2001gat,n1999gat,II3211,n2663gat,n3018gat,n2448gat,n2662gat,
    n2444gat,II3235,n2238gat,n3019gat,n1310gat,n199gat,n87gat,n195gat,n184gat,
    n204gat,II3273,n2168gat,n2452gat,n1691gat,II3287,n3020gat,II3290,n3021gat,
    II3293,n3022gat,n1699gat,II3297,n3023gat,II3300,n3024gat,II3303,n3025gat,
    II3306,n3026gat,II3309,n3027gat,II3312,n3028gat,II3315,n3029gat,II3318,
    n3030gat,n2260gat,n2257gat,n2188gat,n2187gat,n3004gat,II3336,n2039gat,
    II3339,n1774gat,II3342,n1315gat,n2097gat,n1855gat,n2014gat,II3387,n2194gat,
    II3390,n3032gat,n2256gat,II3394,n3033gat,n2251gat,n2184gat,n3003gat,II3401,
    n2192gat,n2133gat,n2131gat,n2185gat,n2049gat,n3001gat,II3412,n2057gat,
    n2253gat,n2252gat,n2248gat,n3006gat,n2264gat,II3429,n2265gat,n2492gat,
    n2329gat,II3436,n1709gat,n1845gat,n1891gat,n1963gat,n1886gat,n1968gat,
    n1958gat,n1629gat,n1895gat,n1631gat,n1711gat,n2990gat,n2200gat,n2078gat,
    n2437gat,n2195gat,II3457,n2556gat,n1956gat,II3461,n3038gat,n1954gat,II3465,
    n3039gat,n1888gat,n2048gat,n2994gat,II3472,n2539gat,n1969gat,n1893gat,
    n1892gat,n2993gat,II3483,n2436gat,n2056gat,n2998gat,II3491,n2387gat,II3494,
    n3043gat,n1960gat,n1887gat,n1961gat,n2996gat,II3504,n2330gat,n2199gat,
    n2147gat,II3509,n3045gat,n2332gat,II3513,n3046gat,n2259gat,n2328gat,
    n3008gat,II3520,n2498gat,n2151gat,n2193gat,n2209gat,n3005gat,II3530,
    n2396gat,n2052gat,n2058gat,n2997gat,II3539,n2198gat,n2349gat,n2215gat,
    n2281gat,n3009gat,II3549,n2197gat,n2146gat,n3002gat,II3558,n2196gat,II3587,
    n2124gat,n2115gat,II3610,n1882gat,II3621,n1974gat,n1955gat,n1970gat,
    n1896gat,n1973gat,n2558gat,n2559gat,II3635,II3646,n2643gat,n2333gat,
    n2564gat,n2352gat,n2642gat,n2636gat,n2637gat,II3660,n88gat,n84gat,n375gat,
    n110gat,II3677,n155gat,n253gat,n1702gat,n150gat,II3691,n151gat,n243gat,
    n233gat,n154gat,n800gat,n2874gat,II3703,n2917gat,n235gat,n2878gat,II3713,
    n2892gat,n372gat,n212gat,n329gat,II3736,n387gat,n334gat,n1700gat,n386gat,
    II3742,n330gat,n1430gat,n1490gat,n452gat,n2885gat,II3754,n2900gat,n333gat,
    n2883gat,II3765,n2929gat,II3777,n462gat,n325gat,n457gat,n2884gat,n461gat,
    n458gat,n2902gat,II3801,n2925gat,n144gat,n247gat,II3808,n326gat,n878gat,
    n2879gat,II3817,n2916gat,n382gat,II3831,n383gat,n134gat,n2875gat,II3841,
    n2899gat,n254gat,n252gat,n2877gat,n468gat,II3867,n469gat,n381gat,n2893gat,
    II3876,n2926gat,n241gat,n140gat,II3882,n255gat,n802gat,n2882gat,II3891,
    n2924gat,n146gat,II3904,n147gat,n380gat,n2881gat,II3914,n2923gat,n69gat,
    n68gat,n1885gat,II3923,n2710gat,n2707gat,n16gat,n295gat,n357gat,n11gat,
    n12gat,n1889gat,II3935,n2704gat,n2700gat,n2051gat,II3941,n2684gat,n2680gat,
    n1350gat,II3945,n2696gat,II3948,n2692gat,II3951,n2683gat,II3954,n2679gat,
    II3957,n2449gat,n1754gat,II3962,n2830gat,n2827gat,n2512gat,n1544gat,
    n1769gat,n1683gat,n1756gat,n2167gat,n2013gat,II4000,n1791gat,n2691gat,
    n2695gat,n1518gat,n2699gat,n2703gat,n2159gat,n2478gat,II4014,n2744gat,
    n2740gat,n2158gat,n2186gat,II4020,n2800gat,n2797gat,n2288gat,II4024,
    n1513gat,n2537gat,n2538gat,n2442gat,n2483gat,n1334gat,II4055,n1747gat,
    II4067,n1674gat,n1403gat,n1402gat,II4081,n1806gat,n1634gat,n1338gat,II4105,
    n1455gat,II4108,n1339gat,n1505gat,n2980gat,II4117,n2758gat,n2755gat,
    n1546gat,II4122,n2752gat,n2748gat,n2012gat,n2016gat,n2002gat,n2008gat,
    II4129,n2858gat,n2857gat,II4135,n2766gat,II4138,n2765gat,n1684gat,n1759gat,
    II4145,II4157,n1524gat,n1862gat,n1863gat,n1919gat,n1860gat,n1460gat,II4185,
    n1595gat,n1454gat,n1469gat,n1468gat,n1519gat,II4194,n1461gat,n1477gat,
    n2984gat,n1594gat,II4212,n1587gat,n1681gat,II4217,II4222,n1761gat,n2751gat,
    n2747gat,II4227,n1760gat,n2743gat,n2739gat,n1978gat,II4233,n1721gat,
    n2808gat,II4236,n2804gat,n517gat,n518gat,n417gat,n418gat,n413gat,n411gat,
    n412gat,n522gat,n406gat,n516gat,n407gat,n355gat,n290gat,n525gat,n527gat,
    n356gat,n416gat,n415gat,n528gat,n521gat,n358gat,n532gat,n639gat,n523gat,
    n1111gat,n635gat,n524gat,n414gat,n1112gat,n630gat,n741gat,n629gat,n633gat,
    n634gat,n926gat,n632gat,n670gat,n636gat,n1123gat,n1007gat,n1006gat,II4309,
    n2941gat,n2814gat,II4312,n2811gat,n1002gat,n2946gat,II4329,n2950gat,
    n2813gat,II4332,n2810gat,n888gat,n2933gat,II4349,n2935gat,n2818gat,II4352,
    n2816gat,n898gat,n2940gat,II4369,n2937gat,n2817gat,II4372,n2815gat,
    n1179gat,n2947gat,II4389,n2956gat,n2824gat,II4392,n2821gat,n897gat,
    n2939gat,II4409,n2938gat,n2823gat,II4412,n2820gat,n894gat,n2932gat,II4429,
    n2936gat,n2829gat,II4432,n2826gat,n1180gat,n2948gat,II4449,n2955gat,
    n2828gat,II4452,n2825gat,n671gat,n628gat,n631gat,n976gat,II4475,n2951gat,
    n2807gat,II4478,n2803gat,n2127gat,II4482,n2682gat,II4485,n2678gat,n2046gat,
    II4489,n2681gat,II4492,n2677gat,n1708gat,II4496,n2688gat,II4499,n2686gat,
    n455gat,n291gat,n2237gat,II4506,n2764gat,n2763gat,n1782gat,II4512,n2762gat,
    n2760gat,n2325gat,II4518,n2761gat,n2759gat,n2245gat,II4524,n2757gat,
    n2754gat,n2244gat,II4530,n2756gat,n2753gat,n2243gat,II4536,n2750gat,
    n2746gat,n2246gat,II4542,n2749gat,n2745gat,n2384gat,II4548,n2742gat,
    n2738gat,n2385gat,II4554,n2741gat,n2737gat,n1286gat,II4558,n2687gat,
    n2685gat,n1328gat,n1381gat,n1384gat,II4566,n2694gat,n2690gat,n1382gat,
    n1451gat,n1453gat,II4573,n2693gat,n2689gat,n927gat,n925gat,n1452gat,II4580,
    n2702gat,n2698gat,n923gat,n921gat,n1890gat,II4587,n2701gat,n2697gat,
    n850gat,n739gat,n1841gat,II4594,n2709gat,n2706gat,n922gat,n848gat,n2047gat,
    II4601,n2708gat,n2705gat,n924gat,n849gat,n2050gat,II4608,n2799gat,n2796gat,
    n1118gat,n1032gat,n2054gat,II4615,n2798gat,n2795gat,II4620,n1745gat,
    n2806gat,II4623,n2802gat,II4626,n1870gat,n1086gat,II4630,n2805gat,II4633,
    n2801gat,n67gat,n85gat,n71gat,n180gat,n1840gat,II4642,n2812gat,n2809gat,
    n76gat,n82gat,n14gat,n186gat,n1842gat,II4651,n2822gat,n2819gat,II4654,
    II4657,II4660,II4663,II4666,II4669,II4672,II4675,II4678,II4681,II4684,
    II4687,II4690,II4693,II4696,II4699,II4702,II4705,II4708,II4711,II4714,
    II4717,II4720,II4723,II4726,II4729,II4732,II4735,II4738,II4741,II4744,
    II4747,II4750,II4753,II4756,II4759,II4762,II4765,II4768,II4771,II4774,
    II4777,II4780,II4783,II4786,II4789,II4792,II4795,II4798,n648gat,n442gat,
    n1214gat,n1215gat,n1216gat,n1217gat,n745gat,n638gat,n423gat,n362gat,
    n749gat,n750gat,n751gat,n752gat,n259gat,n260gat,n261gat,n262gat,n1014gat,
    n1015gat,n1016gat,n1017gat,n476gat,n477gat,n478gat,n479gat,n44gat,n45gat,
    n46gat,n47gat,n168gat,n169gat,n170gat,n171gat,n907gat,n908gat,n909gat,
    n910gat,n344gat,n345gat,n346gat,n347gat,n56gat,n57gat,n58gat,n59gat,
    n768gat,n655gat,n963gat,n868gat,n962gat,n959gat,n945gat,n946gat,n947gat,
    n948gat,n647gat,n441gat,n967gat,n792gat,n1229gat,n1230gat,n1231gat,
    n1232gat,n443gat,n439gat,n966gat,n790gat,n444gat,n440gat,n1051gat,n1052gat,
    n1053gat,n1054gat,n934gat,n935gat,n936gat,n937gat,n710gat,n711gat,n712gat,
    n713gat,n729gat,n730gat,n731gat,n732gat,n494gat,n495gat,n496gat,n497gat,
    n505gat,n506gat,n507gat,n508gat,II1277,n767gat,n653gat,n867gat,n771gat,
    n964gat,n961gat,n804gat,n805gat,n806gat,n807gat,n587gat,n588gat,n589gat,
    n590gat,n447gat,n445gat,n687gat,n688gat,n689gat,n690gat,n568gat,n569gat,
    n570gat,n571gat,II1515,II1584,n1692gat,II1723,II1733,n2428gat,n769gat,
    n1076gat,n766gat,n1185gat,n1186gat,n1187gat,n1188gat,n645gat,n646gat,
    n1383gat,n1327gat,n651gat,n652gat,n765gat,n1202gat,n1203gat,n1204gat,
    n1205gat,n1270gat,n1271gat,n1272gat,n1273gat,n763gat,n1287gat,n1285gat,
    n793gat,n556gat,n795gat,n656gat,n794gat,n773gat,n965gat,n960gat,n780gat,
    n781gat,n782gat,n783gat,n555gat,n450gat,n654gat,n557gat,n874gat,n132gat,
    n649gat,n449gat,n791gat,n650gat,n774gat,n764gat,n222gat,n223gat,n224gat,
    n225gat,n121gat,n122gat,n123gat,n124gat,n2460gat,n2423gat,n2569gat,
    n2570gat,n2571gat,n2572gat,n2410gat,n2411gat,n2412gat,n2413gat,n2580gat,
    n2581gat,n2567gat,n2499gat,n299gat,n207gat,n2647gat,n2648gat,n2602gat,
    n2603gat,n2604gat,n2605gat,n2546gat,n2547gat,n2548gat,n2549gat,n2614gat,
    n2615gat,n2461gat,n2421gat,n2930gat,n1153gat,n1151gat,n982gat,n877gat,
    n2957gat,n1159gat,n1158gat,n1156gat,n1155gat,n1443gat,n1325gat,n1321gat,
    n1320gat,n1368gat,n1258gat,n1373gat,n1372gat,n2978gat,n1441gat,n1440gat,
    n1371gat,n1367gat,n2982gat,n1504gat,n1502gat,n1250gat,n1103gat,n1304gat,
    n1249gat,n1246gat,n1161gat,n1291gat,n1245gat,n2973gat,n1352gat,n1351gat,
    n1303gat,n1302gat,n1163gat,n1102gat,n1101gat,n996gat,n1104gat,n887gat,
    n1305gat,n1162gat,n2977gat,n1360gat,n1359gat,n1358gat,n1357gat,II2720,
    II2735,II2812,n1703gat,n1778gat,n1609gat,II2831,II2889,II2925,II2934,
    n1733gat,n1581gat,n2079gat,n2073gat,n1574gat,n1573gat,n2992gat,n1723gat,
    n1647gat,n1646gat,n2986gat,n1650gat,n1649gat,n1563gat,n2991gat,n1654gat,
    n1653gat,n1644gat,II3148,II3178,n2981gat,n1413gat,n1408gat,n1407gat,
    n2258gat,n2255gat,n2132gat,n2130gat,n3007gat,n2250gat,n2249gat,n1710gat,
    n1630gat,n1894gat,n1847gat,n1846gat,n2055gat,n1967gat,n1959gat,n1957gat,
    n2211gat,n2210gat,n2053gat,n1964gat,n2350gat,n2282gat,n2213gat,n2150gat,
    n2149gat,n2995gat,n1962gat,n2999gat,n1972gat,n1971gat,n3011gat,n2331gat,
    n3015gat,n2566gat,n2565gat,n141gat,n38gat,n37gat,n1074gat,n872gat,n234gat,
    n137gat,n378gat,n377gat,n250gat,n249gat,n248gat,n869gat,n453gat,n448gat,
    n251gat,n244gat,n974gat,n973gat,n870gat,n246gat,n245gat,n460gat,n459gat,
    n975gat,n972gat,n969gat,n145gat,n143gat,n971gat,n970gat,n968gat,n142gat,
    n40gat,n39gat,n772gat,n451gat,n446gat,n139gat,n136gat,n391gat,n390gat,
    n1083gat,n1077gat,n242gat,n240gat,n871gat,n797gat,n324gat,n238gat,n237gat,
    n1082gat,n796gat,n1599gat,II3999,n1586gat,n1755gat,II4023,n1470gat,
    n1400gat,n1399gat,n1398gat,II4144,n1467gat,n1466gat,n2985gat,n1686gat,
    n1533gat,n1532gat,n1531gat,II4216,n2931gat,n1100gat,n994gat,n989gat,
    n880gat,n2943gat,n1012gat,n905gat,n1003gat,n902gat,n1099gat,n998gat,
    n995gat,n980gat,n2960gat,n1175gat,n1174gat,n1001gat,n999gat,n2969gat,
    n1323gat,n1264gat,n981gat,n890gat,n889gat,n886gat,n892gat,n891gat,n2942gat,
    n904gat,n903gat,n1152gat,n1092gat,n997gat,n993gat,n900gat,n895gat,n1094gat,
    n1093gat,n988gat,n984gat,n2965gat,n1267gat,n1257gat,n1178gat,n1116gat,
    n2961gat,n1375gat,n1324gat,n1091gat,n1088gat,n992gat,n987gat,n899gat,
    n896gat,n2967gat,n1262gat,n1260gat,n1098gat,n1090gat,n986gat,n885gat,
    n901gat,n893gat,n1097gat,n1089gat,n1087gat,n991gat,n2968gat,n1326gat,
    n1261gat,n1177gat,n1115gat,n2944gat,n977gat,n2945gat,n1096gat,n1095gat,
    n990gat,n979gat,n2962gat,n1176gat,n1173gat,n1004gat,n1000gat,n1029gat,
    n1028gat,n1031gat,n1030gat,n1011gat,n1181gat,n1010gat,n1005gat,n1182gat,
    n73gat,n70gat,n77gat,n13gat,n1935gat,n197gat,n22gat,n93gat,n2239gat,
    n2433gat,n2427gat,n2583gat,n2650gat,n2617gat,n1598gat,n1154gat,n1411gat,
    n1498gat,n1607gat,n1428gat,n1794gat,n1796gat,n1792gat,n1406gat,n2664gat,
    n1926gat,n1916gat,n1994gat,n1924gat,n1758gat,n200gat,n196gat,n2018gat,
    n89gat,n1471gat,n1472gat,n1600gat,n1397gat,n2005gat,n1818gat,n1510gat,
    n1459gat,n1458gat,n1602gat,n520gat,n519gat,n410gat,n354gat,n408gat,n526gat,
    n531gat,n530gat,n359gat,n420gat,n801gat,n879gat,n1255gat,n1009gat,n409gat,
    n292gat,n419gat,n1243gat,n1171gat,n1244gat,n1265gat,n1254gat,n1008gat,
    n1253gat,n1266gat,n1200gat,n1172gat,n1251gat,n1259gat,n1212gat,n1263gat,
    n978gat,n1199gat,n1252gat,n1757gat;

  dff DFF_0(CK,n673gat,n2897gat);
  dff DFF_1(CK,n398gat,n2782gat);
  dff DFF_2(CK,n402gat,n2790gat);
  dff DFF_3(CK,n919gat,n2670gat);
  dff DFF_4(CK,n846gat,n2793gat);
  dff DFF_5(CK,n394gat,n2782gat);
  dff DFF_6(CK,n703gat,n2790gat);
  dff DFF_7(CK,n722gat,n2670gat);
  dff DFF_8(CK,n726gat,n2793gat);
  dff DFF_9(CK,n2510gat,n748gat);
  dff DFF_10(CK,n271gat,n2732gat);
  dff DFF_11(CK,n160gat,n2776gat);
  dff DFF_12(CK,n337gat,n2735gat);
  dff DFF_13(CK,n842gat,n2673gat);
  dff DFF_14(CK,n341gat,n2779gat);
  dff DFF_15(CK,n2522gat,n43gat);
  dff DFF_16(CK,n2472gat,n1620gat);
  dff DFF_17(CK,n2319gat,n2470gat);
  dff DFF_18(CK,n1821gat,n1827gat);
  dff DFF_19(CK,n1825gat,n1827gat);
  dff DFF_20(CK,n2029gat,n1816gat);
  dff DFF_21(CK,n1829gat,n2027gat);
  dff DFF_22(CK,n283gat,n2732gat);
  dff DFF_23(CK,n165gat,n2776gat);
  dff DFF_24(CK,n279gat,n2735gat);
  dff DFF_25(CK,n1026gat,n2673gat);
  dff DFF_26(CK,n275gat,n2779gat);
  dff DFF_27(CK,n2476gat,n55gat);
  dff DFF_28(CK,n1068gat,n2914gat);
  dff DFF_29(CK,n957gat,n2928gat);
  dff DFF_30(CK,n861gat,n2927gat);
  dff DFF_31(CK,n1294gat,n2896gat);
  dff DFF_32(CK,n1241gat,n2922gat);
  dff DFF_33(CK,n1298gat,n2897gat);
  dff DFF_34(CK,n865gat,n2894gat);
  dff DFF_35(CK,n1080gat,n2921gat);
  dff DFF_36(CK,n1148gat,n2895gat);
  dff DFF_37(CK,n2468gat,n933gat);
  dff DFF_38(CK,n618gat,n2790gat);
  dff DFF_39(CK,n491gat,n2782gat);
  dff DFF_40(CK,n622gat,n2793gat);
  dff DFF_41(CK,n626gat,n2670gat);
  dff DFF_42(CK,n834gat,n3064gat);
  dff DFF_43(CK,n707gat,n3055gat);
  dff DFF_44(CK,n838gat,n3063gat);
  dff DFF_45(CK,n830gat,n3062gat);
  dff DFF_46(CK,n614gat,n3056gat);
  dff DFF_47(CK,n2526gat,n504gat);
  dff DFF_48(CK,n680gat,n2913gat);
  dff DFF_49(CK,n816gat,n2920gat);
  dff DFF_50(CK,n580gat,n2905gat);
  dff DFF_51(CK,n824gat,n3057gat);
  dff DFF_52(CK,n820gat,n3059gat);
  dff DFF_53(CK,n883gat,n3058gat);
  dff DFF_54(CK,n584gat,n2898gat);
  dff DFF_55(CK,n684gat,n3060gat);
  dff DFF_56(CK,n699gat,n3061gat);
  dff DFF_57(CK,n2464gat,n567gat);
  dff DFF_58(CK,n2399gat,n3048gat);
  dff DFF_59(CK,n2343gat,n3049gat);
  dff DFF_60(CK,n2203gat,n3051gat);
  dff DFF_61(CK,n2562gat,n3047gat);
  dff DFF_62(CK,n2207gat,n3050gat);
  dff DFF_63(CK,n2626gat,n3040gat);
  dff DFF_64(CK,n2490gat,n3044gat);
  dff DFF_65(CK,n2622gat,n3042gat);
  dff DFF_66(CK,n2630gat,n3037gat);
  dff DFF_67(CK,n2543gat,n3041gat);
  dff DFF_68(CK,n2102gat,n1606gat);
  dff DFF_69(CK,n1880gat,n3052gat);
  dff DFF_70(CK,n1763gat,n1610gat);
  dff DFF_71(CK,n2155gat,n1858gat);
  dff DFF_72(CK,n1035gat,n2918gat);
  dff DFF_73(CK,n1121gat,n2952gat);
  dff DFF_74(CK,n1072gat,n2919gat);
  dff DFF_75(CK,n1282gat,n2910gat);
  dff DFF_76(CK,n1226gat,n2907gat);
  dff DFF_77(CK,n931gat,n2911gat);
  dff DFF_78(CK,n1135gat,n2912gat);
  dff DFF_79(CK,n1045gat,n2909gat);
  dff DFF_80(CK,n1197gat,n2908gat);
  dff DFF_81(CK,n2518gat,n2971gat);
  dff DFF_82(CK,n667gat,n2904gat);
  dff DFF_83(CK,n659gat,n2891gat);
  dff DFF_84(CK,n553gat,n2903gat);
  dff DFF_85(CK,n777gat,n2915gat);
  dff DFF_86(CK,n561gat,n2901gat);
  dff DFF_87(CK,n366gat,n2890gat);
  dff DFF_88(CK,n322gat,n2888gat);
  dff DFF_89(CK,n318gat,n2887gat);
  dff DFF_90(CK,n314gat,n2886gat);
  dff DFF_91(CK,n2599gat,n3010gat);
  dff DFF_92(CK,n2588gat,n3016gat);
  dff DFF_93(CK,n2640gat,n3054gat);
  dff DFF_94(CK,n2658gat,n2579gat);
  dff DFF_95(CK,n2495gat,n3036gat);
  dff DFF_96(CK,n2390gat,n3034gat);
  dff DFF_97(CK,n2270gat,n3031gat);
  dff DFF_98(CK,n2339gat,n3035gat);
  dff DFF_99(CK,n2502gat,n2646gat);
  dff DFF_100(CK,n2634gat,n3053gat);
  dff DFF_101(CK,n2506gat,n2613gat);
  dff DFF_102(CK,n1834gat,n1625gat);
  dff DFF_103(CK,n1767gat,n1626gat);
  dff DFF_104(CK,n2084gat,n1603gat);
  dff DFF_105(CK,n2143gat,n2541gat);
  dff DFF_106(CK,n2061gat,n2557gat);
  dff DFF_107(CK,n2139gat,n2487gat);
  dff DFF_108(CK,n1899gat,n2532gat);
  dff DFF_109(CK,n1850gat,n2628gat);
  dff DFF_110(CK,n2403gat,n2397gat);
  dff DFF_111(CK,n2394gat,n2341gat);
  dff DFF_112(CK,n2440gat,n2560gat);
  dff DFF_113(CK,n2407gat,n2205gat);
  dff DFF_114(CK,n2347gat,n2201gat);
  dff DFF_115(CK,n1389gat,n1793gat);
  dff DFF_116(CK,n2021gat,n1781gat);
  dff DFF_117(CK,n1394gat,n1516gat);
  dff DFF_118(CK,n1496gat,n1392gat);
  dff DFF_119(CK,n2091gat,n1685gat);
  dff DFF_120(CK,n1332gat,n1565gat);
  dff DFF_121(CK,n1740gat,n1330gat);
  dff DFF_122(CK,n2179gat,n1945gat);
  dff DFF_123(CK,n2190gat,n2268gat);
  dff DFF_124(CK,n2135gat,n2337gat);
  dff DFF_125(CK,n2262gat,n2388gat);
  dff DFF_126(CK,n2182gat,n1836gat);
  dff DFF_127(CK,n1433gat,n2983gat);
  dff DFF_128(CK,n1316gat,n1431gat);
  dff DFF_129(CK,n1363gat,n1314gat);
  dff DFF_130(CK,n1312gat,n1361gat);
  dff DFF_131(CK,n1775gat,n1696gat);
  dff DFF_132(CK,n1871gat,n2009gat);
  dff DFF_133(CK,n2592gat,n1773gat);
  dff DFF_134(CK,n1508gat,n1636gat);
  dff DFF_135(CK,n1678gat,n1712gat);
  dff DFF_136(CK,n2309gat,n3000gat);
  dff DFF_137(CK,n2450gat,n2307gat);
  dff DFF_138(CK,n2446gat,n2661gat);
  dff DFF_139(CK,n2095gat,n827gat);
  dff DFF_140(CK,n2176gat,n2093gat);
  dff DFF_141(CK,n2169gat,n2174gat);
  dff DFF_142(CK,n2454gat,n2163gat);
  dff DFF_143(CK,n2040gat,n1777gat);
  dff DFF_144(CK,n2044gat,n2015gat);
  dff DFF_145(CK,n2037gat,n2042gat);
  dff DFF_146(CK,n2025gat,n2017gat);
  dff DFF_147(CK,n2099gat,n2023gat);
  dff DFF_148(CK,n2266gat,n2493gat);
  dff DFF_149(CK,n2033gat,n2035gat);
  dff DFF_150(CK,n2110gat,n2031gat);
  dff DFF_151(CK,n2125gat,n2108gat);
  dff DFF_152(CK,n2121gat,n2123gat);
  dff DFF_153(CK,n2117gat,n2119gat);
  dff DFF_154(CK,n1975gat,n2632gat);
  dff DFF_155(CK,n2644gat,n2638gat);
  dff DFF_156(CK,n156gat,n612gat);
  dff DFF_157(CK,n152gat,n705gat);
  dff DFF_158(CK,n331gat,n822gat);
  dff DFF_159(CK,n388gat,n881gat);
  dff DFF_160(CK,n463gat,n818gat);
  dff DFF_161(CK,n327gat,n682gat);
  dff DFF_162(CK,n384gat,n697gat);
  dff DFF_163(CK,n256gat,n836gat);
  dff DFF_164(CK,n470gat,n828gat);
  dff DFF_165(CK,n148gat,n832gat);
  dff DFF_166(CK,n2458gat,n2590gat);
  dff DFF_167(CK,n2514gat,n2456gat);
  dff DFF_168(CK,n1771gat,n1613gat);
  dff DFF_169(CK,n1336gat,n1391gat);
  dff DFF_170(CK,n1748gat,n1927gat);
  dff DFF_171(CK,n1675gat,n1713gat);
  dff DFF_172(CK,n1807gat,n1717gat);
  dff DFF_173(CK,n1340gat,n1567gat);
  dff DFF_174(CK,n1456gat,n1564gat);
  dff DFF_175(CK,n1525gat,n1632gat);
  dff DFF_176(CK,n1462gat,n1915gat);
  dff DFF_177(CK,n1596gat,n1800gat);
  dff DFF_178(CK,n1588gat,n1593gat);
assign II1 = ~n3088gat;
assign n2717gat = ~II1;
assign n2715gat = ~n2717gat;
assign II5 = ~n3087gat;
assign n2725gat = ~II5;
assign n2723gat = ~n2725gat;
assign n296gat = ~n421gat;
assign II11 = ~n3093gat;
assign n2768gat = ~II11;
assign II14 = ~n2768gat;
assign n2767gat = ~II14;
assign n373gat = ~n2767gat;
assign II18 = ~n3072gat;
assign n2671gat = ~II18;
assign n2669gat = ~n2671gat;
assign II23 = ~n3081gat;
assign n2845gat = ~II23;
assign n2844gat = ~n2845gat;
assign II27 = ~n3095gat;
assign n2668gat = ~II27;
assign II30 = ~n2668gat;
assign n2667gat = ~II30;
assign n856gat = ~n2667gat;
assign II44 = ~n673gat;
assign n672gat = ~II44;
assign II47 = ~n3069gat;
assign n2783gat = ~II47;
assign II50 = ~n2783gat;
assign n2782gat = ~II50;
assign n396gat = ~n398gat;
assign II62 = ~n3070gat;
assign n2791gat = ~II62;
assign II65 = ~n2791gat;
assign n2790gat = ~II65;
assign II76 = ~n402gat;
assign n401gat = ~II76;
assign n1645gat = ~n1499gat;
assign II81 = ~n2671gat;
assign n2670gat = ~II81;
assign II92 = ~n919gat;
assign n918gat = ~II92;
assign n1553gat = ~n1616gat;
assign II97 = ~n3071gat;
assign n2794gat = ~II97;
assign II100 = ~n2794gat;
assign n2793gat = ~II100;
assign II111 = ~n846gat;
assign n845gat = ~II111;
assign n1559gat = ~n1614gat;
assign n1643gat = ~n1641gat;
assign n1651gat = ~n1642gat;
assign n1562gat = ~n1556gat;
assign n1560gat = ~n1557gat;
assign n1640gat = ~n1639gat;
assign n1566gat = ~n1605gat;
assign n1554gat = ~n1555gat;
assign n1722gat = ~n1558gat;
assign n392gat = ~n394gat;
assign II149 = ~n703gat;
assign n702gat = ~II149;
assign n1319gat = ~n1256gat;
assign n720gat = ~n722gat;
assign II171 = ~n726gat;
assign n725gat = ~II171;
assign n1447gat = ~n1117gat;
assign n1627gat = ~n1618gat;
assign II178 = ~n722gat;
assign n721gat = ~II178;
assign n1380gat = ~n1114gat;
assign n1628gat = ~n1621gat;
assign n701gat = ~n703gat;
assign n1446gat = ~n1318gat;
assign n1705gat = ~n1619gat;
assign n1706gat = ~n1622gat;
assign II192 = ~n3083gat;
assign n2856gat = ~II192;
assign n2854gat = ~n2856gat;
assign II196 = ~n2854gat;
assign n1218gat = ~II196;
assign II199 = ~n3085gat;
assign n2861gat = ~II199;
assign n2859gat = ~n2861gat;
assign II203 = ~n2859gat;
assign n1219gat = ~II203;
assign II206 = ~n3084gat;
assign n2864gat = ~II206;
assign n2862gat = ~n2864gat;
assign II210 = ~n2862gat;
assign n1220gat = ~II210;
assign II214 = ~n2861gat;
assign n2860gat = ~II214;
assign II217 = ~n2860gat;
assign n1221gat = ~II217;
assign II220 = ~n2864gat;
assign n2863gat = ~II220;
assign II223 = ~n2863gat;
assign n1222gat = ~II223;
assign II227 = ~n2856gat;
assign n2855gat = ~II227;
assign II230 = ~n2855gat;
assign n1223gat = ~II230;
assign n640gat = ~n1213gat;
assign II237 = ~n640gat;
assign n753gat = ~II237;
assign II240 = ~n2717gat;
assign n2716gat = ~II240;
assign II243 = ~n3089gat;
assign n2869gat = ~II243;
assign n2867gat = ~n2869gat;
assign II248 = ~n2869gat;
assign n2868gat = ~II248;
assign II253 = ~n2906gat;
assign n754gat = ~II253;
assign II256 = ~n2725gat;
assign n2724gat = ~II256;
assign II259 = ~n3086gat;
assign n2728gat = ~II259;
assign n2726gat = ~n2728gat;
assign II264 = ~n2728gat;
assign n2727gat = ~II264;
assign n422gat = ~n2889gat;
assign II270 = ~n422gat;
assign n755gat = ~II270;
assign n747gat = ~n2906gat;
assign II275 = ~n747gat;
assign n756gat = ~II275;
assign II278 = ~n2889gat;
assign n757gat = ~II278;
assign II282 = ~n1213gat;
assign n758gat = ~II282;
assign n2508gat = ~n2510gat;
assign II297 = ~n3065gat;
assign n2733gat = ~II297;
assign II300 = ~n2733gat;
assign n2732gat = ~II300;
assign II311 = ~n271gat;
assign n270gat = ~II311;
assign II314 = ~n270gat;
assign n263gat = ~II314;
assign II317 = ~n3067gat;
assign n2777gat = ~II317;
assign II320 = ~n2777gat;
assign n2776gat = ~II320;
assign II331 = ~n160gat;
assign n159gat = ~II331;
assign II334 = ~n159gat;
assign n264gat = ~II334;
assign II337 = ~n3066gat;
assign n2736gat = ~II337;
assign II340 = ~n2736gat;
assign n2735gat = ~II340;
assign II351 = ~n337gat;
assign n336gat = ~II351;
assign II354 = ~n336gat;
assign n265gat = ~II354;
assign n158gat = ~n160gat;
assign II359 = ~n158gat;
assign n266gat = ~II359;
assign n335gat = ~n337gat;
assign II363 = ~n335gat;
assign n267gat = ~II363;
assign n269gat = ~n271gat;
assign II368 = ~n269gat;
assign n268gat = ~II368;
assign n41gat = ~n258gat;
assign II375 = ~n41gat;
assign n48gat = ~II375;
assign II378 = ~n725gat;
assign n1018gat = ~II378;
assign II381 = ~n3073gat;
assign n2674gat = ~II381;
assign II384 = ~n2674gat;
assign n2673gat = ~II384;
assign II395 = ~n842gat;
assign n841gat = ~II395;
assign II398 = ~n841gat;
assign n1019gat = ~II398;
assign II401 = ~n721gat;
assign n1020gat = ~II401;
assign n840gat = ~n842gat;
assign II406 = ~n840gat;
assign n1021gat = ~II406;
assign II409 = ~n720gat;
assign n1022gat = ~II409;
assign n724gat = ~n726gat;
assign II414 = ~n724gat;
assign n1023gat = ~II414;
assign II420 = ~n1013gat;
assign n49gat = ~II420;
assign II423 = ~n3068gat;
assign n2780gat = ~II423;
assign II426 = ~n2780gat;
assign n2779gat = ~II426;
assign II437 = ~n341gat;
assign n340gat = ~II437;
assign II440 = ~n340gat;
assign n480gat = ~II440;
assign II443 = ~n702gat;
assign n481gat = ~II443;
assign II446 = ~n394gat;
assign n393gat = ~II446;
assign II449 = ~n393gat;
assign n482gat = ~II449;
assign II453 = ~n701gat;
assign n483gat = ~II453;
assign II456 = ~n392gat;
assign n484gat = ~II456;
assign n339gat = ~n341gat;
assign II461 = ~n339gat;
assign n485gat = ~II461;
assign n42gat = ~n475gat;
assign II468 = ~n42gat;
assign n50gat = ~II468;
assign n162gat = ~n1013gat;
assign II473 = ~n162gat;
assign n51gat = ~II473;
assign II476 = ~n475gat;
assign n52gat = ~II476;
assign II480 = ~n258gat;
assign n53gat = ~II480;
assign n2520gat = ~n2522gat;
assign n1448gat = ~n1376gat;
assign n1701gat = ~n1617gat;
assign n1379gat = ~n1377gat;
assign n1615gat = ~n1624gat;
assign n1500gat = ~n1113gat;
assign n1503gat = ~n1501gat;
assign n1779gat = ~n1623gat;
assign II509 = ~n3099gat;
assign n2730gat = ~II509;
assign II512 = ~n2730gat;
assign n2729gat = ~II512;
assign n2470gat = ~n2472gat;
assign n2317gat = ~n2319gat;
assign n1819gat = ~n1821gat;
assign n1823gat = ~n1825gat;
assign n1816gat = ~n1817gat;
assign n2027gat = ~n2029gat;
assign II572 = ~n1829gat;
assign n1828gat = ~II572;
assign II576 = ~n3100gat;
assign n2851gat = ~II576;
assign II579 = ~n2851gat;
assign n2850gat = ~II579;
assign II583 = ~n2786gat;
assign n2785gat = ~II583;
assign n92gat = ~n2785gat;
assign n637gat = ~n529gat;
assign n293gat = ~n361gat;
assign II591 = ~n3094gat;
assign n2722gat = ~II591;
assign II594 = ~n2722gat;
assign n2721gat = ~II594;
assign n297gat = ~n2721gat;
assign II606 = ~n283gat;
assign n282gat = ~II606;
assign II609 = ~n282gat;
assign n172gat = ~II609;
assign II620 = ~n165gat;
assign n164gat = ~II620;
assign II623 = ~n164gat;
assign n173gat = ~II623;
assign II634 = ~n279gat;
assign n278gat = ~II634;
assign II637 = ~n278gat;
assign n174gat = ~II637;
assign n163gat = ~n165gat;
assign II642 = ~n163gat;
assign n175gat = ~II642;
assign n277gat = ~n279gat;
assign II646 = ~n277gat;
assign n176gat = ~II646;
assign n281gat = ~n283gat;
assign II651 = ~n281gat;
assign n177gat = ~II651;
assign n54gat = ~n167gat;
assign II658 = ~n54gat;
assign n60gat = ~II658;
assign II661 = ~n845gat;
assign n911gat = ~II661;
assign II672 = ~n1026gat;
assign n1025gat = ~II672;
assign II675 = ~n1025gat;
assign n912gat = ~II675;
assign II678 = ~n918gat;
assign n913gat = ~II678;
assign n1024gat = ~n1026gat;
assign II683 = ~n1024gat;
assign n914gat = ~II683;
assign n917gat = ~n919gat;
assign II687 = ~n917gat;
assign n915gat = ~II687;
assign n844gat = ~n846gat;
assign II692 = ~n844gat;
assign n916gat = ~II692;
assign II698 = ~n906gat;
assign n61gat = ~II698;
assign II709 = ~n275gat;
assign n274gat = ~II709;
assign II712 = ~n274gat;
assign n348gat = ~II712;
assign II715 = ~n401gat;
assign n349gat = ~II715;
assign II718 = ~n398gat;
assign n397gat = ~II718;
assign II721 = ~n397gat;
assign n350gat = ~II721;
assign n400gat = ~n402gat;
assign II726 = ~n400gat;
assign n351gat = ~II726;
assign II729 = ~n396gat;
assign n352gat = ~II729;
assign n273gat = ~n275gat;
assign II734 = ~n273gat;
assign n353gat = ~II734;
assign n178gat = ~n343gat;
assign II741 = ~n178gat;
assign n62gat = ~II741;
assign n66gat = ~n906gat;
assign II746 = ~n66gat;
assign n63gat = ~II746;
assign II749 = ~n343gat;
assign n64gat = ~II749;
assign II753 = ~n167gat;
assign n65gat = ~II753;
assign n2474gat = ~n2476gat;
assign II768 = ~n3090gat;
assign n2832gat = ~II768;
assign II771 = ~n2832gat;
assign n2831gat = ~II771;
assign n2731gat = ~n2733gat;
assign II776 = ~n3074gat;
assign n2719gat = ~II776;
assign n2718gat = ~n2719gat;
assign II790 = ~n1068gat;
assign n1067gat = ~II790;
assign II793 = ~n1067gat;
assign n949gat = ~II793;
assign II796 = ~n3076gat;
assign n2839gat = ~II796;
assign n2838gat = ~n2839gat;
assign n2775gat = ~n2777gat;
assign II812 = ~n957gat;
assign n956gat = ~II812;
assign II815 = ~n956gat;
assign n950gat = ~II815;
assign II818 = ~n3075gat;
assign n2712gat = ~II818;
assign n2711gat = ~n2712gat;
assign n2734gat = ~n2736gat;
assign II834 = ~n861gat;
assign n860gat = ~II834;
assign II837 = ~n860gat;
assign n951gat = ~II837;
assign n955gat = ~n957gat;
assign II842 = ~n955gat;
assign n952gat = ~II842;
assign n859gat = ~n861gat;
assign II846 = ~n859gat;
assign n953gat = ~II846;
assign n1066gat = ~n1068gat;
assign II851 = ~n1066gat;
assign n954gat = ~II851;
assign n857gat = ~n944gat;
assign II858 = ~n857gat;
assign n938gat = ~II858;
assign n2792gat = ~n2794gat;
assign II863 = ~n3080gat;
assign n2847gat = ~II863;
assign n2846gat = ~n2847gat;
assign II877 = ~n1294gat;
assign n1293gat = ~II877;
assign II880 = ~n1293gat;
assign n1233gat = ~II880;
assign n2672gat = ~n2674gat;
assign II885 = ~n3082gat;
assign n2853gat = ~II885;
assign n2852gat = ~n2853gat;
assign II899 = ~n1241gat;
assign n1240gat = ~II899;
assign II902 = ~n1240gat;
assign n1234gat = ~II902;
assign II913 = ~n1298gat;
assign n1297gat = ~II913;
assign II916 = ~n1297gat;
assign n1235gat = ~II916;
assign n1239gat = ~n1241gat;
assign II921 = ~n1239gat;
assign n1236gat = ~II921;
assign n1296gat = ~n1298gat;
assign II925 = ~n1296gat;
assign n1237gat = ~II925;
assign n1292gat = ~n1294gat;
assign II930 = ~n1292gat;
assign n1238gat = ~II930;
assign II936 = ~n1228gat;
assign n939gat = ~II936;
assign n2778gat = ~n2780gat;
assign II941 = ~n3077gat;
assign n2837gat = ~II941;
assign n2836gat = ~n2837gat;
assign II955 = ~n865gat;
assign n864gat = ~II955;
assign II958 = ~n864gat;
assign n1055gat = ~II958;
assign n2789gat = ~n2791gat;
assign II963 = ~n3079gat;
assign n2841gat = ~II963;
assign n2840gat = ~n2841gat;
assign II977 = ~n1080gat;
assign n1079gat = ~II977;
assign II980 = ~n1079gat;
assign n1056gat = ~II980;
assign n2781gat = ~n2783gat;
assign II985 = ~n3078gat;
assign n2843gat = ~II985;
assign n2842gat = ~n2843gat;
assign II999 = ~n1148gat;
assign n1147gat = ~II999;
assign II1002 = ~n1147gat;
assign n1057gat = ~II1002;
assign n1078gat = ~n1080gat;
assign II1007 = ~n1078gat;
assign n1058gat = ~II1007;
assign n1146gat = ~n1148gat;
assign II1011 = ~n1146gat;
assign n1059gat = ~II1011;
assign n863gat = ~n865gat;
assign II1016 = ~n863gat;
assign n1060gat = ~II1016;
assign n928gat = ~n1050gat;
assign II1023 = ~n928gat;
assign n940gat = ~II1023;
assign n858gat = ~n1228gat;
assign II1028 = ~n858gat;
assign n941gat = ~II1028;
assign II1031 = ~n1050gat;
assign n942gat = ~II1031;
assign II1035 = ~n944gat;
assign n943gat = ~II1035;
assign n2466gat = ~n2468gat;
assign n2720gat = ~n2722gat;
assign n740gat = ~n2667gat;
assign n2784gat = ~n2786gat;
assign n743gat = ~n746gat;
assign n294gat = ~n360gat;
assign n374gat = ~n2767gat;
assign n616gat = ~n618gat;
assign II1067 = ~n616gat;
assign n501gat = ~II1067;
assign n489gat = ~n491gat;
assign II1079 = ~n489gat;
assign n502gat = ~II1079;
assign II1082 = ~n618gat;
assign n617gat = ~II1082;
assign II1085 = ~n617gat;
assign n499gat = ~II1085;
assign II1088 = ~n491gat;
assign n490gat = ~II1088;
assign II1091 = ~n490gat;
assign n500gat = ~II1091;
assign n620gat = ~n622gat;
assign II1103 = ~n620gat;
assign n738gat = ~II1103;
assign n624gat = ~n626gat;
assign II1115 = ~n624gat;
assign n737gat = ~II1115;
assign II1118 = ~n622gat;
assign n621gat = ~II1118;
assign II1121 = ~n621gat;
assign n733gat = ~II1121;
assign II1124 = ~n626gat;
assign n625gat = ~II1124;
assign II1127 = ~n625gat;
assign n735gat = ~II1127;
assign II1138 = ~n834gat;
assign n833gat = ~II1138;
assign II1141 = ~n833gat;
assign n714gat = ~II1141;
assign II1152 = ~n707gat;
assign n706gat = ~II1152;
assign II1155 = ~n706gat;
assign n715gat = ~II1155;
assign II1166 = ~n838gat;
assign n837gat = ~II1166;
assign II1169 = ~n837gat;
assign n716gat = ~II1169;
assign n705gat = ~n707gat;
assign II1174 = ~n705gat;
assign n717gat = ~II1174;
assign n836gat = ~n838gat;
assign II1178 = ~n836gat;
assign n718gat = ~II1178;
assign n832gat = ~n834gat;
assign II1183 = ~n832gat;
assign n719gat = ~II1183;
assign n515gat = ~n709gat;
assign II1190 = ~n515gat;
assign n509gat = ~II1190;
assign II1201 = ~n830gat;
assign n829gat = ~II1201;
assign II1204 = ~n829gat;
assign n734gat = ~II1204;
assign n828gat = ~n830gat;
assign II1209 = ~n828gat;
assign n736gat = ~II1209;
assign II1216 = ~n728gat;
assign n510gat = ~II1216;
assign II1227 = ~n614gat;
assign n613gat = ~II1227;
assign II1230 = ~n613gat;
assign n498gat = ~II1230;
assign n612gat = ~n614gat;
assign II1236 = ~n612gat;
assign n503gat = ~II1236;
assign n404gat = ~n493gat;
assign II1243 = ~n404gat;
assign n511gat = ~II1243;
assign n405gat = ~n728gat;
assign II1248 = ~n405gat;
assign n512gat = ~II1248;
assign II1251 = ~n493gat;
assign n513gat = ~II1251;
assign II1255 = ~n709gat;
assign n514gat = ~II1255;
assign n2524gat = ~n2526gat;
assign n17gat = ~n564gat;
assign n79gat = ~n86gat;
assign n219gat = ~n78gat;
assign n563gat = ~II1278;
assign n289gat = ~n563gat;
assign n179gat = ~n287gat;
assign n188gat = ~n288gat;
assign n72gat = ~n181gat;
assign n111gat = ~n182gat;
assign II1302 = ~n680gat;
assign n679gat = ~II1302;
assign II1305 = ~n679gat;
assign n808gat = ~II1305;
assign II1319 = ~n816gat;
assign n815gat = ~II1319;
assign II1322 = ~n815gat;
assign n809gat = ~II1322;
assign II1336 = ~n580gat;
assign n579gat = ~II1336;
assign II1339 = ~n579gat;
assign n810gat = ~II1339;
assign n814gat = ~n816gat;
assign II1344 = ~n814gat;
assign n811gat = ~II1344;
assign n578gat = ~n580gat;
assign II1348 = ~n578gat;
assign n812gat = ~II1348;
assign n678gat = ~n680gat;
assign II1353 = ~n678gat;
assign n813gat = ~II1353;
assign n677gat = ~n803gat;
assign II1360 = ~n677gat;
assign n572gat = ~II1360;
assign II1371 = ~n824gat;
assign n823gat = ~II1371;
assign II1374 = ~n823gat;
assign n591gat = ~II1374;
assign II1385 = ~n820gat;
assign n819gat = ~II1385;
assign II1388 = ~n819gat;
assign n592gat = ~II1388;
assign II1399 = ~n883gat;
assign n882gat = ~II1399;
assign II1402 = ~n882gat;
assign n593gat = ~II1402;
assign n818gat = ~n820gat;
assign II1407 = ~n818gat;
assign n594gat = ~II1407;
assign n881gat = ~n883gat;
assign II1411 = ~n881gat;
assign n595gat = ~II1411;
assign n822gat = ~n824gat;
assign II1416 = ~n822gat;
assign n596gat = ~II1416;
assign II1422 = ~n586gat;
assign n573gat = ~II1422;
assign II1436 = ~n584gat;
assign n583gat = ~II1436;
assign II1439 = ~n583gat;
assign n691gat = ~II1439;
assign II1450 = ~n684gat;
assign n683gat = ~II1450;
assign II1453 = ~n683gat;
assign n692gat = ~II1453;
assign II1464 = ~n699gat;
assign n698gat = ~II1464;
assign II1467 = ~n698gat;
assign n693gat = ~II1467;
assign n682gat = ~n684gat;
assign II1472 = ~n682gat;
assign n694gat = ~II1472;
assign n697gat = ~n699gat;
assign II1476 = ~n697gat;
assign n695gat = ~II1476;
assign n582gat = ~n584gat;
assign II1481 = ~n582gat;
assign n696gat = ~II1481;
assign n456gat = ~n686gat;
assign II1488 = ~n456gat;
assign n574gat = ~II1488;
assign n565gat = ~n586gat;
assign II1493 = ~n565gat;
assign n575gat = ~II1493;
assign II1496 = ~n686gat;
assign n576gat = ~II1496;
assign II1500 = ~n803gat;
assign n577gat = ~II1500;
assign n2462gat = ~n2464gat;
assign n2665gat = ~II1516;
assign n2596gat = ~n2665gat;
assign n189gat = ~n286gat;
assign n194gat = ~n187gat;
assign n21gat = ~n15gat;
assign II1538 = ~n2399gat;
assign n2398gat = ~II1538;
assign n2353gat = ~n2398gat;
assign II1550 = ~n2343gat;
assign n2342gat = ~II1550;
assign n2284gat = ~n2342gat;
assign n2201gat = ~n2203gat;
assign n2354gat = ~n2201gat;
assign n2560gat = ~n2562gat;
assign n2356gat = ~n2560gat;
assign n2205gat = ~n2207gat;
assign n2214gat = ~n2205gat;
assign n2286gat = ~II1585;
assign n2624gat = ~n2626gat;
assign II1606 = ~n2490gat;
assign n2489gat = ~II1606;
assign II1617 = ~n2622gat;
assign n2621gat = ~II1617;
assign n2533gat = ~n2534gat;
assign II1630 = ~n2630gat;
assign n2629gat = ~II1630;
assign n2486gat = ~n2629gat;
assign n2541gat = ~n2543gat;
assign n2429gat = ~n2541gat;
assign n2432gat = ~n2430gat;
assign II1655 = ~n2102gat;
assign n2101gat = ~II1655;
assign n1693gat = ~n2101gat;
assign II1667 = ~n1880gat;
assign n1879gat = ~II1667;
assign n1698gat = ~n1934gat;
assign n1543gat = ~n1606gat;
assign II1683 = ~n1763gat;
assign n1762gat = ~II1683;
assign n1673gat = ~n2989gat;
assign n1858gat = ~n1673gat;
assign II1698 = ~n2155gat;
assign n2154gat = ~II1698;
assign n2488gat = ~n2490gat;
assign II1703 = ~n2626gat;
assign n2625gat = ~II1703;
assign n2530gat = ~n2531gat;
assign II1708 = ~n2543gat;
assign n2542gat = ~II1708;
assign n2482gat = ~n2542gat;
assign n2426gat = ~n2480gat;
assign n2153gat = ~n2155gat;
assign n2341gat = ~n2343gat;
assign n2355gat = ~n2341gat;
assign II1719 = ~n2562gat;
assign n2561gat = ~II1719;
assign n2443gat = ~n2561gat;
assign n2289gat = ~II1724;
assign n2148gat = ~II1734;
assign n855gat = ~n2148gat;
assign n759gat = ~n855gat;
assign II1749 = ~n1035gat;
assign n1034gat = ~II1749;
assign II1752 = ~n1034gat;
assign n1189gat = ~II1752;
assign n1075gat = ~n855gat;
assign II1766 = ~n1121gat;
assign n1120gat = ~II1766;
assign II1769 = ~n1120gat;
assign n1190gat = ~II1769;
assign n760gat = ~n855gat;
assign II1783 = ~n1072gat;
assign n1071gat = ~II1783;
assign II1786 = ~n1071gat;
assign n1191gat = ~II1786;
assign n1119gat = ~n1121gat;
assign II1791 = ~n1119gat;
assign n1192gat = ~II1791;
assign n1070gat = ~n1072gat;
assign II1795 = ~n1070gat;
assign n1193gat = ~II1795;
assign n1033gat = ~n1035gat;
assign II1800 = ~n1033gat;
assign n1194gat = ~II1800;
assign n1183gat = ~n1184gat;
assign II1807 = ~n1183gat;
assign n1274gat = ~II1807;
assign n644gat = ~n855gat;
assign n1280gat = ~n1282gat;
assign n641gat = ~n855gat;
assign II1833 = ~n1226gat;
assign n1225gat = ~II1833;
assign II1837 = ~n1282gat;
assign n1281gat = ~II1837;
assign n1224gat = ~n1226gat;
assign II1843 = ~n2970gat;
assign n1275gat = ~II1843;
assign n761gat = ~n855gat;
assign II1857 = ~n931gat;
assign n930gat = ~II1857;
assign II1860 = ~n930gat;
assign n1206gat = ~II1860;
assign n762gat = ~n855gat;
assign II1874 = ~n1135gat;
assign n1134gat = ~II1874;
assign II1877 = ~n1134gat;
assign n1207gat = ~II1877;
assign n643gat = ~n855gat;
assign II1891 = ~n1045gat;
assign n1044gat = ~II1891;
assign II1894 = ~n1044gat;
assign n1208gat = ~II1894;
assign n1133gat = ~n1135gat;
assign II1899 = ~n1133gat;
assign n1209gat = ~II1899;
assign n1043gat = ~n1045gat;
assign II1903 = ~n1043gat;
assign n1210gat = ~II1903;
assign n929gat = ~n931gat;
assign II1908 = ~n929gat;
assign n1211gat = ~II1908;
assign n1268gat = ~n1201gat;
assign II1915 = ~n1268gat;
assign n1276gat = ~II1915;
assign n1329gat = ~n2970gat;
assign II1920 = ~n1329gat;
assign n1277gat = ~II1920;
assign II1923 = ~n1201gat;
assign n1278gat = ~II1923;
assign II1927 = ~n1184gat;
assign n1279gat = ~II1927;
assign n1284gat = ~n1269gat;
assign n642gat = ~n855gat;
assign n1195gat = ~n1197gat;
assign II1947 = ~n1197gat;
assign n1196gat = ~II1947;
assign n2516gat = ~n2518gat;
assign II1961 = ~n2516gat;
assign n3017gat = ~II1961;
assign n851gat = ~n853gat;
assign n1725gat = ~n2148gat;
assign n664gat = ~n1725gat;
assign n852gat = ~n854gat;
assign II1981 = ~n667gat;
assign n666gat = ~II1981;
assign n368gat = ~n1725gat;
assign II1996 = ~n659gat;
assign n658gat = ~II1996;
assign II1999 = ~n658gat;
assign n784gat = ~II1999;
assign n662gat = ~n1725gat;
assign II2014 = ~n553gat;
assign n552gat = ~II2014;
assign II2017 = ~n552gat;
assign n785gat = ~II2017;
assign n661gat = ~n1725gat;
assign II2032 = ~n777gat;
assign n776gat = ~II2032;
assign II2035 = ~n776gat;
assign n786gat = ~II2035;
assign n551gat = ~n553gat;
assign II2040 = ~n551gat;
assign n787gat = ~II2040;
assign n775gat = ~n777gat;
assign II2044 = ~n775gat;
assign n788gat = ~II2044;
assign n657gat = ~n659gat;
assign II2049 = ~n657gat;
assign n789gat = ~II2049;
assign n35gat = ~n779gat;
assign II2056 = ~n35gat;
assign n125gat = ~II2056;
assign n558gat = ~n1725gat;
assign n559gat = ~n561gat;
assign n371gat = ~n1725gat;
assign II2084 = ~n366gat;
assign n365gat = ~II2084;
assign II2088 = ~n561gat;
assign n560gat = ~II2088;
assign n364gat = ~n366gat;
assign II2094 = ~n2876gat;
assign n126gat = ~II2094;
assign n663gat = ~n1725gat;
assign II2109 = ~n322gat;
assign n321gat = ~II2109;
assign II2112 = ~n321gat;
assign n226gat = ~II2112;
assign n370gat = ~n1725gat;
assign II2127 = ~n318gat;
assign n317gat = ~II2127;
assign II2130 = ~n317gat;
assign n227gat = ~II2130;
assign n369gat = ~n1725gat;
assign II2145 = ~n314gat;
assign n313gat = ~II2145;
assign II2148 = ~n313gat;
assign n228gat = ~II2148;
assign n316gat = ~n318gat;
assign II2153 = ~n316gat;
assign n229gat = ~II2153;
assign n312gat = ~n314gat;
assign II2157 = ~n312gat;
assign n230gat = ~II2157;
assign n320gat = ~n322gat;
assign II2162 = ~n320gat;
assign n231gat = ~II2162;
assign n34gat = ~n221gat;
assign II2169 = ~n34gat;
assign n127gat = ~II2169;
assign n133gat = ~n2876gat;
assign II2174 = ~n133gat;
assign n128gat = ~II2174;
assign II2177 = ~n221gat;
assign n129gat = ~II2177;
assign II2181 = ~n779gat;
assign n130gat = ~II2181;
assign n665gat = ~n667gat;
assign n1601gat = ~n120gat;
assign n2597gat = ~n2599gat;
assign n2595gat = ~n2594gat;
assign n2586gat = ~n2588gat;
assign II2213 = ~n2342gat;
assign n2573gat = ~II2213;
assign n2638gat = ~n2640gat;
assign II2225 = ~n2638gat;
assign n2574gat = ~II2225;
assign II2228 = ~n2561gat;
assign n2575gat = ~II2228;
assign II2232 = ~n2640gat;
assign n2639gat = ~II2232;
assign II2235 = ~n2639gat;
assign n2576gat = ~II2235;
assign II2238 = ~n2560gat;
assign n2577gat = ~II2238;
assign II2242 = ~n2341gat;
assign n2578gat = ~II2242;
assign II2248 = ~n2568gat;
assign n2582gat = ~II2248;
assign II2251 = ~n2207gat;
assign n2206gat = ~II2251;
assign II2254 = ~n2206gat;
assign n2414gat = ~II2254;
assign II2257 = ~n2398gat;
assign n2415gat = ~II2257;
assign II2260 = ~n2203gat;
assign n2202gat = ~II2260;
assign II2263 = ~n2202gat;
assign n2416gat = ~II2263;
assign n2397gat = ~n2399gat;
assign II2268 = ~n2397gat;
assign n2417gat = ~II2268;
assign II2271 = ~n2201gat;
assign n2418gat = ~II2271;
assign II2275 = ~n2205gat;
assign n2419gat = ~II2275;
assign II2281 = ~n2409gat;
assign n2585gat = ~II2281;
assign n2656gat = ~n2658gat;
assign n2493gat = ~n2495gat;
assign n2388gat = ~n2390gat;
assign II2316 = ~n2390gat;
assign n2389gat = ~II2316;
assign II2319 = ~n2495gat;
assign n2494gat = ~II2319;
assign II2324 = ~n3014gat;
assign n2649gat = ~II2324;
assign n2268gat = ~n2270gat;
assign II2344 = ~n2339gat;
assign n2338gat = ~II2344;
assign n2337gat = ~n2339gat;
assign II2349 = ~n2270gat;
assign n2269gat = ~II2349;
assign II2354 = ~n2880gat;
assign n2652gat = ~II2354;
assign n2500gat = ~n2502gat;
assign n2620gat = ~n2622gat;
assign n2612gat = ~n2620gat;
assign II2372 = ~n2612gat;
assign n2606gat = ~II2372;
assign n2532gat = ~n2625gat;
assign II2376 = ~n2532gat;
assign n2607gat = ~II2376;
assign n2540gat = ~n2488gat;
assign II2380 = ~n2540gat;
assign n2608gat = ~II2380;
assign n2536gat = ~n2624gat;
assign II2385 = ~n2536gat;
assign n2609gat = ~II2385;
assign n2487gat = ~n2489gat;
assign II2389 = ~n2487gat;
assign n2610gat = ~II2389;
assign n2557gat = ~n2621gat;
assign II2394 = ~n2557gat;
assign n2611gat = ~II2394;
assign II2400 = ~n2601gat;
assign n2616gat = ~II2400;
assign II2403 = ~n2629gat;
assign n2550gat = ~II2403;
assign II2414 = ~n2634gat;
assign n2633gat = ~II2414;
assign II2417 = ~n2633gat;
assign n2551gat = ~II2417;
assign II2420 = ~n2542gat;
assign n2552gat = ~II2420;
assign n2632gat = ~n2634gat;
assign II2425 = ~n2632gat;
assign n2553gat = ~II2425;
assign II2428 = ~n2541gat;
assign n2554gat = ~II2428;
assign n2628gat = ~n2630gat;
assign II2433 = ~n2628gat;
assign n2555gat = ~II2433;
assign II2439 = ~n2545gat;
assign n2619gat = ~II2439;
assign n2504gat = ~n2506gat;
assign n2660gat = ~n2655gat;
assign n1528gat = ~n2293gat;
assign n1523gat = ~n2219gat;
assign n1592gat = ~n1529gat;
assign n2666gat = ~n1704gat;
assign n2422gat = ~n3013gat;
assign n2290gat = ~n2202gat;
assign n2081gat = ~n2218gat;
assign n2285gat = ~n2397gat;
assign n2359gat = ~n2358gat;
assign n1414gat = ~n1415gat;
assign n566gat = ~n364gat;
assign n1480gat = ~n2292gat;
assign n1301gat = ~n1416gat;
assign n1150gat = ~n312gat;
assign n873gat = ~n316gat;
assign n2011gat = ~n2306gat;
assign n1478gat = ~n1481gat;
assign n875gat = ~n559gat;
assign n1410gat = ~n2357gat;
assign n876gat = ~n1347gat;
assign n1160gat = ~n1484gat;
assign n1084gat = ~n657gat;
assign n983gat = ~n320gat;
assign n1482gat = ~n2363gat;
assign n1157gat = ~n1483gat;
assign n985gat = ~n775gat;
assign n1530gat = ~n2364gat;
assign n1307gat = ~n1308gat;
assign n1085gat = ~n551gat;
assign n1479gat = ~n2291gat;
assign n1348gat = ~n1349gat;
assign n2217gat = ~n2206gat;
assign n1591gat = ~n2223gat;
assign n1437gat = ~n1438gat;
assign n1832gat = ~n1834gat;
assign n1765gat = ~n1767gat;
assign n1878gat = ~n1880gat;
assign n1442gat = ~n1831gat;
assign n1444gat = ~n1442gat;
assign n1378gat = ~n2975gat;
assign n1322gat = ~n2974gat;
assign n1439gat = ~n1486gat;
assign n1370gat = ~n1426gat;
assign n1369gat = ~n2966gat;
assign n1366gat = ~n1365gat;
assign n1374gat = ~n2979gat;
assign n2162gat = ~n2220gat;
assign n1450gat = ~n1423gat;
assign n1427gat = ~n1608gat;
assign n1603gat = ~n1831gat;
assign n2082gat = ~n2084gat;
assign n1449gat = ~n1494gat;
assign n1590gat = ~n1603gat;
assign n1248gat = ~n2954gat;
assign n1418gat = ~n1417gat;
assign n1306gat = ~n2964gat;
assign n1353gat = ~n1419gat;
assign n1247gat = ~n2958gat;
assign n1355gat = ~n1422gat;
assign n1300gat = ~n2963gat;
assign n1487gat = ~n1485gat;
assign n1164gat = ~n2953gat;
assign n1356gat = ~n1354gat;
assign n1436gat = ~n1435gat;
assign n1106gat = ~n2949gat;
assign n1425gat = ~n1421gat;
assign n1105gat = ~n2934gat;
assign n1424gat = ~n1420gat;
assign n1309gat = ~n2959gat;
assign II2672 = ~n2143gat;
assign n2142gat = ~II2672;
assign n1788gat = ~n2142gat;
assign II2684 = ~n2061gat;
assign n2060gat = ~II2684;
assign n1786gat = ~n2060gat;
assign II2696 = ~n2139gat;
assign n2138gat = ~II2696;
assign n1839gat = ~n2138gat;
assign n1897gat = ~n1899gat;
assign n1884gat = ~n1897gat;
assign n1848gat = ~n1850gat;
assign n1783gat = ~n1848gat;
assign n1548gat = ~II2721;
assign n1719gat = ~n1548gat;
assign n2137gat = ~n2139gat;
assign n1633gat = ~n2137gat;
assign n2059gat = ~n2061gat;
assign n1785gat = ~n2059gat;
assign II2731 = ~n1850gat;
assign n1849gat = ~II2731;
assign n1784gat = ~n1849gat;
assign n1716gat = ~II2736;
assign n1635gat = ~n1716gat;
assign n2401gat = ~n2403gat;
assign n1989gat = ~n2401gat;
assign n2392gat = ~n2394gat;
assign n1918gat = ~n2392gat;
assign II2771 = ~n2440gat;
assign n2439gat = ~II2771;
assign n1986gat = ~n2439gat;
assign n1866gat = ~n1865gat;
assign II2785 = ~n2407gat;
assign n2406gat = ~II2785;
assign n2216gat = ~n2406gat;
assign n2345gat = ~n2347gat;
assign n1988gat = ~n2345gat;
assign n1735gat = ~n1861gat;
assign n1387gat = ~n1389gat;
assign n1694gat = ~II2813;
assign n1777gat = ~n1694gat;
assign n1781gat = ~n1780gat;
assign n2019gat = ~n2021gat;
assign n1549gat = ~II2832;
assign n1551gat = ~n1549gat;
assign II2837 = ~n2347gat;
assign n2346gat = ~II2837;
assign n2152gat = ~n2346gat;
assign n2405gat = ~n2407gat;
assign n2351gat = ~n2405gat;
assign II2843 = ~n2403gat;
assign n2402gat = ~II2843;
assign n2212gat = ~n2402gat;
assign II2847 = ~n2394gat;
assign n2393gat = ~II2847;
assign n1991gat = ~n2393gat;
assign n1665gat = ~n1666gat;
assign n1517gat = ~n1578gat;
assign n1392gat = ~n1394gat;
assign II2873 = ~n1496gat;
assign n1495gat = ~II2873;
assign n1685gat = ~n1604gat;
assign II2885 = ~n2091gat;
assign n2090gat = ~II2885;
assign n1550gat = ~II2890;
assign n1552gat = ~n1550gat;
assign n1330gat = ~n1332gat;
assign n1738gat = ~n1740gat;
assign II2915 = ~n1740gat;
assign n1739gat = ~II2915;
assign n1925gat = ~n1920gat;
assign n1917gat = ~n1921gat;
assign n2141gat = ~n2143gat;
assign n1787gat = ~n2141gat;
assign n1717gat = ~II2926;
assign n1859gat = ~n1717gat;
assign n1922gat = ~n1798gat;
assign n1713gat = ~II2935;
assign n1743gat = ~n1713gat;
assign n1923gat = ~n1864gat;
assign n1945gat = ~n1690gat;
assign II2953 = ~n2179gat;
assign n2178gat = ~II2953;
assign n1661gat = ~n1660gat;
assign n1572gat = ~n1576gat;
assign n2438gat = ~n2440gat;
assign n2283gat = ~n2438gat;
assign n1520gat = ~n1582gat;
assign n1580gat = ~n1577gat;
assign n1990gat = ~n2988gat;
assign II2978 = ~n2190gat;
assign n2189gat = ~II2978;
assign II2989 = ~n2135gat;
assign n2134gat = ~II2989;
assign II3000 = ~n2262gat;
assign n2261gat = ~II3000;
assign n2128gat = ~n2129gat;
assign n1836gat = ~n1695gat;
assign II3016 = ~n2182gat;
assign n2181gat = ~II3016;
assign n1431gat = ~n1433gat;
assign n1314gat = ~n1316gat;
assign n1361gat = ~n1363gat;
assign II3056 = ~n1312gat;
assign n1311gat = ~II3056;
assign n1707gat = ~n1626gat;
assign n1773gat = ~n1775gat;
assign n1659gat = ~n2987gat;
assign n1515gat = ~n1521gat;
assign n1736gat = ~n1737gat;
assign n1658gat = ~n2216gat;
assign n1724gat = ~n1732gat;
assign n1662gat = ~n1663gat;
assign n1656gat = ~n1655gat;
assign n1670gat = ~n1667gat;
assign n1569gat = ~n1570gat;
assign n1568gat = ~n1575gat;
assign n1727gat = ~n1728gat;
assign n1797gat = ~n1801gat;
assign n1730gat = ~n1731gat;
assign n1561gat = ~n1571gat;
assign n1668gat = ~n1734gat;
assign n1742gat = ~n2216gat;
assign n1671gat = ~n1669gat;
assign n1652gat = ~n1657gat;
assign n1648gat = ~n1729gat;
assign n1790gat = ~n1726gat;
assign n2004gat = ~n1929gat;
assign n1869gat = ~n1871gat;
assign II3143 = ~n2592gat;
assign n2591gat = ~II3143;
assign n1584gat = ~n2989gat;
assign n1714gat = ~II3149;
assign n1718gat = ~n1714gat;
assign II3163 = ~n1508gat;
assign n1507gat = ~II3163;
assign n1396gat = ~n1401gat;
assign II3168 = ~n1394gat;
assign n1393gat = ~II3168;
assign n1409gat = ~n1476gat;
assign II3174 = ~n1899gat;
assign n1898gat = ~II3174;
assign n1838gat = ~n1898gat;
assign n1712gat = ~II3179;
assign II3191 = ~n1678gat;
assign n1677gat = ~II3191;
assign n2000gat = ~n1412gat;
assign n2001gat = ~n1412gat;
assign n1999gat = ~n2001gat;
assign n2307gat = ~n2309gat;
assign II3211 = ~n2663gat;
assign n3018gat = ~II3211;
assign n2448gat = ~n2450gat;
assign n2661gat = ~n2662gat;
assign n2444gat = ~n2446gat;
assign II3235 = ~n2238gat;
assign n3019gat = ~II3235;
assign n1310gat = ~n1312gat;
assign n199gat = ~n87gat;
assign n195gat = ~n184gat;
assign n827gat = ~n204gat;
assign n2093gat = ~n2095gat;
assign n2174gat = ~n2176gat;
assign II3273 = ~n2169gat;
assign n2168gat = ~II3273;
assign n2452gat = ~n2454gat;
assign n1691gat = ~n2452gat;
assign II3287 = ~n1691gat;
assign n3020gat = ~II3287;
assign II3290 = ~n1691gat;
assign n3021gat = ~II3290;
assign II3293 = ~n1691gat;
assign n3022gat = ~II3293;
assign n1699gat = ~n2452gat;
assign II3297 = ~n1699gat;
assign n3023gat = ~II3297;
assign II3300 = ~n1699gat;
assign n3024gat = ~II3300;
assign II3303 = ~n1691gat;
assign n3025gat = ~II3303;
assign II3306 = ~n1699gat;
assign n3026gat = ~II3306;
assign II3309 = ~n1699gat;
assign n3027gat = ~II3309;
assign II3312 = ~n1699gat;
assign n3028gat = ~II3312;
assign II3315 = ~n1869gat;
assign n3029gat = ~II3315;
assign II3318 = ~n1869gat;
assign n3030gat = ~II3318;
assign n2260gat = ~n2262gat;
assign n2257gat = ~n2189gat;
assign n2188gat = ~n2190gat;
assign n2187gat = ~n3004gat;
assign II3336 = ~n2040gat;
assign n2039gat = ~II3336;
assign II3339 = ~n1775gat;
assign n1774gat = ~II3339;
assign II3342 = ~n1316gat;
assign n1315gat = ~II3342;
assign n2042gat = ~n2044gat;
assign n2035gat = ~n2037gat;
assign n2023gat = ~n2025gat;
assign n2097gat = ~n2099gat;
assign n1855gat = ~n2014gat;
assign II3387 = ~n2194gat;
assign n3031gat = ~II3387;
assign II3390 = ~n2261gat;
assign n3032gat = ~II3390;
assign n2256gat = ~n3032gat;
assign II3394 = ~n2260gat;
assign n3033gat = ~II3394;
assign n2251gat = ~n3033gat;
assign n2184gat = ~n3003gat;
assign II3401 = ~n2192gat;
assign n3034gat = ~II3401;
assign n2133gat = ~n2135gat;
assign n2131gat = ~n2185gat;
assign n2049gat = ~n3001gat;
assign II3412 = ~n2057gat;
assign n3035gat = ~II3412;
assign n2253gat = ~n2189gat;
assign n2252gat = ~n2260gat;
assign n2248gat = ~n3006gat;
assign n2264gat = ~n2266gat;
assign II3429 = ~n2266gat;
assign n2265gat = ~II3429;
assign n2492gat = ~n2329gat;
assign II3436 = ~n2492gat;
assign n3036gat = ~II3436;
assign n1709gat = ~n1849gat;
assign n1845gat = ~n2141gat;
assign n1891gat = ~n2059gat;
assign n1963gat = ~n2137gat;
assign n1886gat = ~n1897gat;
assign n1968gat = ~n1958gat;
assign n1629gat = ~n1895gat;
assign n1631gat = ~n1848gat;
assign n1711gat = ~n2990gat;
assign n2200gat = ~n2078gat;
assign n2437gat = ~n2195gat;
assign II3457 = ~n2556gat;
assign n3037gat = ~II3457;
assign n1956gat = ~n1898gat;
assign II3461 = ~n1956gat;
assign n3038gat = ~II3461;
assign n1954gat = ~n3038gat;
assign II3465 = ~n1886gat;
assign n3039gat = ~II3465;
assign n1888gat = ~n3039gat;
assign n2048gat = ~n2994gat;
assign II3472 = ~n2539gat;
assign n3040gat = ~II3472;
assign n1969gat = ~n2142gat;
assign n1893gat = ~n2060gat;
assign n1892gat = ~n2993gat;
assign II3483 = ~n2436gat;
assign n3041gat = ~II3483;
assign n2056gat = ~n2998gat;
assign II3491 = ~n2387gat;
assign n3042gat = ~II3491;
assign II3494 = ~n1963gat;
assign n3043gat = ~II3494;
assign n1960gat = ~n3043gat;
assign n1887gat = ~n2138gat;
assign n1961gat = ~n2996gat;
assign II3504 = ~n2330gat;
assign n3044gat = ~II3504;
assign n2199gat = ~n2147gat;
assign II3509 = ~n2438gat;
assign n3045gat = ~II3509;
assign n2332gat = ~n3045gat;
assign II3513 = ~n2439gat;
assign n3046gat = ~II3513;
assign n2259gat = ~n3046gat;
assign n2328gat = ~n3008gat;
assign II3520 = ~n2498gat;
assign n3047gat = ~II3520;
assign n2151gat = ~n2193gat;
assign n2209gat = ~n3005gat;
assign II3530 = ~n2396gat;
assign n3048gat = ~II3530;
assign n2052gat = ~n2393gat;
assign n2058gat = ~n2997gat;
assign II3539 = ~n2198gat;
assign n3049gat = ~II3539;
assign n2349gat = ~n2215gat;
assign n2281gat = ~n3009gat;
assign II3549 = ~n2197gat;
assign n3050gat = ~II3549;
assign n2146gat = ~n3002gat;
assign II3558 = ~n2196gat;
assign n3051gat = ~II3558;
assign n2031gat = ~n2033gat;
assign n2108gat = ~n2110gat;
assign II3587 = ~n2125gat;
assign n2124gat = ~II3587;
assign n2123gat = ~n2125gat;
assign n2119gat = ~n2121gat;
assign n2115gat = ~n2117gat;
assign II3610 = ~n1882gat;
assign n3052gat = ~II3610;
assign II3621 = ~n1975gat;
assign n1974gat = ~II3621;
assign n1955gat = ~n1956gat;
assign n1970gat = ~n1896gat;
assign n1973gat = ~n1975gat;
assign n2558gat = ~n2559gat;
assign II3635 = ~n2558gat;
assign n3053gat = ~II3635;
assign II3646 = ~n2644gat;
assign n2643gat = ~II3646;
assign n2333gat = ~n2438gat;
assign n2564gat = ~n2352gat;
assign n2642gat = ~n2644gat;
assign n2636gat = ~n2637gat;
assign II3660 = ~n2636gat;
assign n3054gat = ~II3660;
assign n88gat = ~n84gat;
assign n375gat = ~n110gat;
assign II3677 = ~n156gat;
assign n155gat = ~II3677;
assign n253gat = ~n1702gat;
assign n150gat = ~n152gat;
assign II3691 = ~n152gat;
assign n151gat = ~II3691;
assign n243gat = ~n1702gat;
assign n233gat = ~n243gat;
assign n154gat = ~n156gat;
assign n800gat = ~n2874gat;
assign II3703 = ~n2917gat;
assign n3055gat = ~II3703;
assign n235gat = ~n2878gat;
assign II3713 = ~n2892gat;
assign n3056gat = ~II3713;
assign n372gat = ~n212gat;
assign n329gat = ~n331gat;
assign II3736 = ~n388gat;
assign n387gat = ~II3736;
assign n334gat = ~n1700gat;
assign n386gat = ~n388gat;
assign II3742 = ~n331gat;
assign n330gat = ~II3742;
assign n1430gat = ~n1700gat;
assign n1490gat = ~n1430gat;
assign n452gat = ~n2885gat;
assign II3754 = ~n2900gat;
assign n3057gat = ~II3754;
assign n333gat = ~n2883gat;
assign II3765 = ~n2929gat;
assign n3058gat = ~II3765;
assign II3777 = ~n463gat;
assign n462gat = ~II3777;
assign n325gat = ~n327gat;
assign n457gat = ~n2884gat;
assign n461gat = ~n463gat;
assign n458gat = ~n2902gat;
assign II3801 = ~n2925gat;
assign n3059gat = ~II3801;
assign n144gat = ~n247gat;
assign II3808 = ~n327gat;
assign n326gat = ~II3808;
assign n878gat = ~n2879gat;
assign II3817 = ~n2916gat;
assign n3060gat = ~II3817;
assign n382gat = ~n384gat;
assign II3831 = ~n384gat;
assign n383gat = ~II3831;
assign n134gat = ~n2875gat;
assign II3841 = ~n2899gat;
assign n3061gat = ~II3841;
assign n254gat = ~n256gat;
assign n252gat = ~n2877gat;
assign n468gat = ~n470gat;
assign II3867 = ~n470gat;
assign n469gat = ~II3867;
assign n381gat = ~n2893gat;
assign II3876 = ~n2926gat;
assign n3062gat = ~II3876;
assign n241gat = ~n140gat;
assign II3882 = ~n256gat;
assign n255gat = ~II3882;
assign n802gat = ~n2882gat;
assign II3891 = ~n2924gat;
assign n3063gat = ~II3891;
assign n146gat = ~n148gat;
assign II3904 = ~n148gat;
assign n147gat = ~II3904;
assign n380gat = ~n2881gat;
assign II3914 = ~n2923gat;
assign n3064gat = ~II3914;
assign n69gat = ~n68gat;
assign n1885gat = ~n2048gat;
assign II3923 = ~n2710gat;
assign n2707gat = ~II3923;
assign n16gat = ~n564gat;
assign n295gat = ~n357gat;
assign n11gat = ~n12gat;
assign n1889gat = ~n1961gat;
assign II3935 = ~n2704gat;
assign n2700gat = ~II3935;
assign n2051gat = ~n2056gat;
assign II3941 = ~n2684gat;
assign n2680gat = ~II3941;
assign n1350gat = ~n1831gat;
assign II3945 = ~n1350gat;
assign n2696gat = ~II3945;
assign II3948 = ~n2696gat;
assign n2692gat = ~II3948;
assign II3951 = ~n2448gat;
assign n2683gat = ~II3951;
assign II3954 = ~n2683gat;
assign n2679gat = ~II3954;
assign II3957 = ~n2450gat;
assign n2449gat = ~II3957;
assign n1754gat = ~n2449gat;
assign II3962 = ~n2830gat;
assign n2827gat = ~II3962;
assign n2590gat = ~n2592gat;
assign n2456gat = ~n2458gat;
assign n2512gat = ~n2514gat;
assign n1544gat = ~n1625gat;
assign n1769gat = ~n1771gat;
assign n1683gat = ~n1756gat;
assign n2167gat = ~n2169gat;
assign n2013gat = ~II4000;
assign n1791gat = ~n2013gat;
assign n2691gat = ~n2695gat;
assign n1518gat = ~n1694gat;
assign n2699gat = ~n2703gat;
assign n2159gat = ~n1412gat;
assign n2478gat = ~n2579gat;
assign II4014 = ~n2744gat;
assign n2740gat = ~II4014;
assign n2158gat = ~n1412gat;
assign n2186gat = ~n2613gat;
assign II4020 = ~n2800gat;
assign n2797gat = ~II4020;
assign n2288gat = ~II4024;
assign n1513gat = ~n2288gat;
assign n2537gat = ~n2538gat;
assign n2442gat = ~n2483gat;
assign n1334gat = ~n1336gat;
assign II4055 = ~n1748gat;
assign n1747gat = ~II4055;
assign II4067 = ~n1675gat;
assign n1674gat = ~II4067;
assign n1403gat = ~n1402gat;
assign II4081 = ~n1807gat;
assign n1806gat = ~II4081;
assign n1634gat = ~n1712gat;
assign n1338gat = ~n1340gat;
assign II4105 = ~n1456gat;
assign n1455gat = ~II4105;
assign II4108 = ~n1340gat;
assign n1339gat = ~II4108;
assign n1505gat = ~n2980gat;
assign II4117 = ~n1505gat;
assign n2758gat = ~II4117;
assign n2755gat = ~n2758gat;
assign n1546gat = ~n2980gat;
assign II4122 = ~n1546gat;
assign n2752gat = ~II4122;
assign n2748gat = ~n2752gat;
assign n2012gat = ~n2016gat;
assign n2002gat = ~n2008gat;
assign II4129 = ~n3097gat;
assign n2858gat = ~II4129;
assign n2857gat = ~n2858gat;
assign II4135 = ~n3098gat;
assign n2766gat = ~II4135;
assign II4138 = ~n2766gat;
assign n2765gat = ~II4138;
assign n1684gat = ~n1759gat;
assign n1632gat = ~II4145;
assign II4157 = ~n1525gat;
assign n1524gat = ~II4157;
assign n1862gat = ~n1863gat;
assign n1919gat = ~n1860gat;
assign n1460gat = ~n1462gat;
assign II4185 = ~n1596gat;
assign n1595gat = ~II4185;
assign n1454gat = ~n1469gat;
assign n1468gat = ~n1519gat;
assign II4194 = ~n1462gat;
assign n1461gat = ~II4194;
assign n1477gat = ~n2984gat;
assign n1594gat = ~n1596gat;
assign II4212 = ~n1588gat;
assign n1587gat = ~II4212;
assign n1681gat = ~II4217;
assign II4222 = ~n1761gat;
assign n2751gat = ~II4222;
assign n2747gat = ~n2751gat;
assign II4227 = ~n1760gat;
assign n2743gat = ~II4227;
assign n2739gat = ~n2743gat;
assign n1978gat = ~n2286gat;
assign II4233 = ~n1721gat;
assign n2808gat = ~II4233;
assign II4236 = ~n2808gat;
assign n2804gat = ~II4236;
assign n517gat = ~n518gat;
assign n417gat = ~n418gat;
assign n413gat = ~n411gat;
assign n412gat = ~n522gat;
assign n406gat = ~n516gat;
assign n407gat = ~n355gat;
assign n290gat = ~n525gat;
assign n527gat = ~n356gat;
assign n416gat = ~n415gat;
assign n528gat = ~n521gat;
assign n358gat = ~n532gat;
assign n639gat = ~n523gat;
assign n1111gat = ~n635gat;
assign n524gat = ~n414gat;
assign n1112gat = ~n630gat;
assign n741gat = ~n629gat;
assign n633gat = ~n634gat;
assign n926gat = ~n632gat;
assign n670gat = ~n636gat;
assign n1123gat = ~n632gat;
assign n1007gat = ~n635gat;
assign n1006gat = ~n630gat;
assign II4309 = ~n2941gat;
assign n2814gat = ~II4309;
assign II4312 = ~n2814gat;
assign n2811gat = ~II4312;
assign n1002gat = ~n2946gat;
assign II4329 = ~n2950gat;
assign n2813gat = ~II4329;
assign II4332 = ~n2813gat;
assign n2810gat = ~II4332;
assign n888gat = ~n2933gat;
assign II4349 = ~n2935gat;
assign n2818gat = ~II4349;
assign II4352 = ~n2818gat;
assign n2816gat = ~II4352;
assign n898gat = ~n2940gat;
assign II4369 = ~n2937gat;
assign n2817gat = ~II4369;
assign II4372 = ~n2817gat;
assign n2815gat = ~II4372;
assign n1179gat = ~n2947gat;
assign II4389 = ~n2956gat;
assign n2824gat = ~II4389;
assign II4392 = ~n2824gat;
assign n2821gat = ~II4392;
assign n897gat = ~n2939gat;
assign II4409 = ~n2938gat;
assign n2823gat = ~II4409;
assign II4412 = ~n2823gat;
assign n2820gat = ~II4412;
assign n894gat = ~n2932gat;
assign II4429 = ~n2936gat;
assign n2829gat = ~II4429;
assign II4432 = ~n2829gat;
assign n2826gat = ~II4432;
assign n1180gat = ~n2948gat;
assign II4449 = ~n2955gat;
assign n2828gat = ~II4449;
assign II4452 = ~n2828gat;
assign n2825gat = ~II4452;
assign n671gat = ~n673gat;
assign n628gat = ~n631gat;
assign n976gat = ~n628gat;
assign II4475 = ~n2951gat;
assign n2807gat = ~II4475;
assign II4478 = ~n2807gat;
assign n2803gat = ~II4478;
assign n2127gat = ~n2389gat;
assign II4482 = ~n2127gat;
assign n2682gat = ~II4482;
assign II4485 = ~n2682gat;
assign n2678gat = ~II4485;
assign n2046gat = ~n2269gat;
assign II4489 = ~n2046gat;
assign n2681gat = ~II4489;
assign II4492 = ~n2681gat;
assign n2677gat = ~II4492;
assign n1708gat = ~n2338gat;
assign II4496 = ~n1708gat;
assign n2688gat = ~II4496;
assign II4499 = ~n2688gat;
assign n2686gat = ~II4499;
assign n455gat = ~n291gat;
assign n2237gat = ~n2646gat;
assign II4506 = ~n2764gat;
assign n2763gat = ~II4506;
assign n1782gat = ~n2971gat;
assign II4512 = ~n2762gat;
assign n2760gat = ~II4512;
assign n2325gat = ~n3010gat;
assign II4518 = ~n2761gat;
assign n2759gat = ~II4518;
assign n2245gat = ~n504gat;
assign II4524 = ~n2757gat;
assign n2754gat = ~II4524;
assign n2244gat = ~n567gat;
assign II4530 = ~n2756gat;
assign n2753gat = ~II4530;
assign n2243gat = ~n55gat;
assign II4536 = ~n2750gat;
assign n2746gat = ~II4536;
assign n2246gat = ~n933gat;
assign II4542 = ~n2749gat;
assign n2745gat = ~II4542;
assign n2384gat = ~n43gat;
assign II4548 = ~n2742gat;
assign n2738gat = ~II4548;
assign n2385gat = ~n748gat;
assign II4554 = ~n2741gat;
assign n2737gat = ~II4554;
assign n1286gat = ~n1269gat;
assign II4558 = ~n1286gat;
assign n2687gat = ~II4558;
assign n2685gat = ~n2687gat;
assign n1328gat = ~n1224gat;
assign n1381gat = ~n1328gat;
assign n1384gat = ~n2184gat;
assign II4566 = ~n2694gat;
assign n2690gat = ~II4566;
assign n1382gat = ~n1280gat;
assign n1451gat = ~n1382gat;
assign n1453gat = ~n2187gat;
assign II4573 = ~n2693gat;
assign n2689gat = ~II4573;
assign n927gat = ~n1133gat;
assign n925gat = ~n927gat;
assign n1452gat = ~n2049gat;
assign II4580 = ~n2702gat;
assign n2698gat = ~II4580;
assign n923gat = ~n1043gat;
assign n921gat = ~n923gat;
assign n1890gat = ~n2328gat;
assign II4587 = ~n2701gat;
assign n2697gat = ~II4587;
assign n850gat = ~n929gat;
assign n739gat = ~n850gat;
assign n1841gat = ~n2058gat;
assign II4594 = ~n2709gat;
assign n2706gat = ~II4594;
assign n922gat = ~n1119gat;
assign n848gat = ~n922gat;
assign n2047gat = ~n2209gat;
assign II4601 = ~n2708gat;
assign n2705gat = ~II4601;
assign n924gat = ~n1070gat;
assign n849gat = ~n924gat;
assign n2050gat = ~n2146gat;
assign II4608 = ~n2799gat;
assign n2796gat = ~II4608;
assign n1118gat = ~n1033gat;
assign n1032gat = ~n1118gat;
assign n2054gat = ~n2281gat;
assign II4615 = ~n2798gat;
assign n2795gat = ~II4615;
assign II4620 = ~n1745gat;
assign n2806gat = ~II4620;
assign II4623 = ~n2806gat;
assign n2802gat = ~II4623;
assign II4626 = ~n1871gat;
assign n1870gat = ~II4626;
assign n1086gat = ~n1870gat;
assign II4630 = ~n1086gat;
assign n2805gat = ~II4630;
assign II4633 = ~n2805gat;
assign n2801gat = ~II4633;
assign n67gat = ~n85gat;
assign n71gat = ~n180gat;
assign n1840gat = ~n1892gat;
assign II4642 = ~n2812gat;
assign n2809gat = ~II4642;
assign n76gat = ~n82gat;
assign n14gat = ~n186gat;
assign n1842gat = ~n1711gat;
assign II4651 = ~n2822gat;
assign n2819gat = ~II4651;
assign II4654 = ~n2819gat;
assign n3104gat = ~II4654;
assign II4657 = ~n2809gat;
assign n3105gat = ~II4657;
assign II4660 = ~n2801gat;
assign n3106gat = ~II4660;
assign II4663 = ~n2802gat;
assign n3107gat = ~II4663;
assign II4666 = ~n2795gat;
assign n3108gat = ~II4666;
assign II4669 = ~n2796gat;
assign n3109gat = ~II4669;
assign II4672 = ~n2705gat;
assign n3110gat = ~II4672;
assign II4675 = ~n2706gat;
assign n3111gat = ~II4675;
assign II4678 = ~n2697gat;
assign n3112gat = ~II4678;
assign II4681 = ~n2698gat;
assign n3113gat = ~II4681;
assign II4684 = ~n2689gat;
assign n3114gat = ~II4684;
assign II4687 = ~n2690gat;
assign n3115gat = ~II4687;
assign II4690 = ~n2685gat;
assign n3116gat = ~II4690;
assign II4693 = ~n2737gat;
assign n3117gat = ~II4693;
assign II4696 = ~n2738gat;
assign n3118gat = ~II4696;
assign II4699 = ~n2745gat;
assign n3119gat = ~II4699;
assign II4702 = ~n2746gat;
assign n3120gat = ~II4702;
assign II4705 = ~n2753gat;
assign n3121gat = ~II4705;
assign II4708 = ~n2754gat;
assign n3122gat = ~II4708;
assign II4711 = ~n2759gat;
assign n3123gat = ~II4711;
assign II4714 = ~n2760gat;
assign n3124gat = ~II4714;
assign II4717 = ~n2763gat;
assign n3125gat = ~II4717;
assign II4720 = ~n2686gat;
assign n3126gat = ~II4720;
assign II4723 = ~n2677gat;
assign n3127gat = ~II4723;
assign II4726 = ~n2678gat;
assign n3128gat = ~II4726;
assign II4729 = ~n2803gat;
assign n3129gat = ~II4729;
assign II4732 = ~n2825gat;
assign n3130gat = ~II4732;
assign II4735 = ~n2826gat;
assign n3131gat = ~II4735;
assign II4738 = ~n2820gat;
assign n3132gat = ~II4738;
assign II4741 = ~n2821gat;
assign n3133gat = ~II4741;
assign II4744 = ~n2815gat;
assign n3134gat = ~II4744;
assign II4747 = ~n2816gat;
assign n3135gat = ~II4747;
assign II4750 = ~n2810gat;
assign n3136gat = ~II4750;
assign II4753 = ~n2811gat;
assign n3137gat = ~II4753;
assign II4756 = ~n2804gat;
assign n3138gat = ~II4756;
assign II4759 = ~n2739gat;
assign n3139gat = ~II4759;
assign II4762 = ~n2747gat;
assign n3140gat = ~II4762;
assign II4765 = ~n2748gat;
assign n3141gat = ~II4765;
assign II4768 = ~n2755gat;
assign n3142gat = ~II4768;
assign II4771 = ~n2797gat;
assign n3143gat = ~II4771;
assign II4774 = ~n2740gat;
assign n3144gat = ~II4774;
assign II4777 = ~n2699gat;
assign n3145gat = ~II4777;
assign II4780 = ~n2691gat;
assign n3146gat = ~II4780;
assign II4783 = ~n2827gat;
assign n3147gat = ~II4783;
assign II4786 = ~n2679gat;
assign n3148gat = ~II4786;
assign II4789 = ~n2692gat;
assign n3149gat = ~II4789;
assign II4792 = ~n2680gat;
assign n3150gat = ~II4792;
assign II4795 = ~n2700gat;
assign n3151gat = ~II4795;
assign II4798 = ~n2707gat;
assign n3152gat = ~II4798;
assign n2897gat = n648gat | n442gat;
assign n1213gat = n1214gat | n1215gat | n1216gat | n1217gat;
assign n2906gat = n745gat | n638gat;
assign n2889gat = n423gat | n362gat;
assign n748gat = n749gat | n750gat | n751gat | n752gat;
assign n258gat = n259gat | n260gat | n261gat | n262gat;
assign n1013gat = n1014gat | n1015gat | n1016gat | n1017gat;
assign n475gat = n476gat | n477gat | n478gat | n479gat;
assign n43gat = n44gat | n45gat | n46gat | n47gat;
assign n2786gat = n3091gat | n3092gat;
assign n167gat = n168gat | n169gat | n170gat | n171gat;
assign n906gat = n907gat | n908gat | n909gat | n910gat;
assign n343gat = n344gat | n345gat | n346gat | n347gat;
assign n55gat = n56gat | n57gat | n58gat | n59gat;
assign n2914gat = n768gat | n655gat;
assign n2928gat = n963gat | n868gat;
assign n2927gat = n962gat | n959gat;
assign n944gat = n945gat | n946gat | n947gat | n948gat;
assign n2896gat = n647gat | n441gat;
assign n2922gat = n967gat | n792gat;
assign n1228gat = n1229gat | n1230gat | n1231gat | n1232gat;
assign n2894gat = n443gat | n439gat;
assign n2921gat = n966gat | n790gat;
assign n2895gat = n444gat | n440gat;
assign n1050gat = n1051gat | n1052gat | n1053gat | n1054gat;
assign n933gat = n934gat | n935gat | n936gat | n937gat;
assign n709gat = n710gat | n711gat | n712gat | n713gat;
assign n728gat = n729gat | n730gat | n731gat | n732gat;
assign n493gat = n494gat | n495gat | n496gat | n497gat;
assign n504gat = n505gat | n506gat | n507gat | n508gat;
assign II1277 = n2860gat | n2855gat | n2863gat;
assign II1278 = n740gat | n3030gat | II1277;
assign n2913gat = n767gat | n653gat;
assign n2920gat = n867gat | n771gat;
assign n2905gat = n964gat | n961gat;
assign n803gat = n804gat | n805gat | n806gat | n807gat;
assign n586gat = n587gat | n588gat | n589gat | n590gat;
assign n2898gat = n447gat | n445gat;
assign n686gat = n687gat | n688gat | n689gat | n690gat;
assign n567gat = n568gat | n569gat | n570gat | n571gat;
assign II1515 = n2474gat | n2524gat | n2831gat;
assign II1516 = n2466gat | n2462gat | II1515;
assign II1584 = n2353gat | n2284gat | n2354gat;
assign II1585 = n2356gat | n2214gat | II1584;
assign n2989gat = n1693gat | n1692gat;
assign II1723 = n2354gat | n2353gat | n2214gat;
assign II1724 = n2355gat | n2443gat | II1723;
assign II1733 = n2286gat | n2428gat | n2289gat;
assign II1734 = n1604gat | n2214gat | II1733;
assign n2918gat = n769gat | n759gat;
assign n2952gat = n1076gat | n1075gat;
assign n2919gat = n766gat | n760gat;
assign n1184gat = n1185gat | n1186gat | n1187gat | n1188gat;
assign n2910gat = n645gat | n644gat;
assign n2907gat = n646gat | n641gat;
assign n2970gat = n1383gat | n1327gat;
assign n2911gat = n761gat | n651gat;
assign n2912gat = n762gat | n652gat;
assign n2909gat = n765gat | n643gat;
assign n1201gat = n1202gat | n1203gat | n1204gat | n1205gat;
assign n1269gat = n1270gat | n1271gat | n1272gat | n1273gat;
assign n2908gat = n763gat | n642gat;
assign n2971gat = n1287gat | n1285gat;
assign n2904gat = n793gat | n664gat | n556gat;
assign n2891gat = n795gat | n656gat | n368gat;
assign n2903gat = n794gat | n773gat | n662gat;
assign n2915gat = n965gat | n960gat | n661gat;
assign n779gat = n780gat | n781gat | n782gat | n783gat;
assign n2901gat = n558gat | n555gat | n450gat;
assign n2890gat = n654gat | n557gat | n371gat;
assign n2876gat = n874gat | n132gat;
assign n2888gat = n663gat | n649gat | n449gat;
assign n2887gat = n791gat | n650gat | n370gat;
assign n2886gat = n774gat | n764gat | n369gat;
assign n221gat = n222gat | n223gat | n224gat | n225gat;
assign n120gat = n121gat | n122gat | n123gat | n124gat;
assign n3010gat = n2460gat | n2423gat;
assign n3016gat = n2596gat | n2595gat;
assign n2568gat = n2569gat | n2570gat | n2571gat | n2572gat;
assign n2409gat = n2410gat | n2411gat | n2412gat | n2413gat;
assign n2579gat = n2580gat | n2581gat;
assign n3014gat = n2567gat | n2499gat;
assign n2880gat = n299gat | n207gat;
assign n2646gat = n2647gat | n2648gat;
assign n2601gat = n2602gat | n2603gat | n2604gat | n2605gat;
assign n2545gat = n2546gat | n2547gat | n2548gat | n2549gat;
assign n2613gat = n2614gat | n2615gat;
assign n3013gat = n2461gat | n2421gat;
assign n2930gat = n1153gat | n1151gat | n982gat | n877gat;
assign n2957gat = n1159gat | n1158gat | n1156gat | n1155gat;
assign n2975gat = n1443gat | n1325gat;
assign n2974gat = n1321gat | n1320gat;
assign n2966gat = n1368gat | n1258gat;
assign n2979gat = n1373gat | n1372gat;
assign n2978gat = n1441gat | n1440gat | n1371gat | n1367gat;
assign n2982gat = n1504gat | n1502gat;
assign n2954gat = n1250gat | n1103gat;
assign n2964gat = n1304gat | n1249gat;
assign n2958gat = n1246gat | n1161gat;
assign n2963gat = n1291gat | n1245gat;
assign n2973gat = n1352gat | n1351gat | n1303gat | n1302gat;
assign n2953gat = n1163gat | n1102gat;
assign n2949gat = n1101gat | n996gat;
assign n2934gat = n1104gat | n887gat;
assign n2959gat = n1305gat | n1162gat;
assign n2977gat = n1360gat | n1359gat | n1358gat | n1357gat;
assign II2720 = n1788gat | n1786gat | n1839gat;
assign II2721 = n1884gat | n1783gat | II2720;
assign II2735 = n1788gat | n1884gat | n1633gat;
assign II2736 = n1785gat | n1784gat | II2735;
assign II2812 = n1703gat | n1704gat | n1778gat;
assign II2813 = n1609gat | n1702gat | n1700gat | II2812;
assign II2831 = n1839gat | n1786gat | n1788gat;
assign II2832 = n1884gat | n1784gat | II2831;
assign II2889 = n1784gat | n1633gat | n1884gat;
assign II2890 = n1788gat | n1786gat | II2889;
assign II2925 = n1784gat | n1785gat | n1633gat;
assign II2926 = n1884gat | n1787gat | II2925;
assign II2934 = n1784gat | n1839gat | n1788gat;
assign II2935 = n1785gat | n1884gat | II2934;
assign n2988gat = n1733gat | n1581gat;
assign n2983gat = n2079gat | n2073gat;
assign n2987gat = n1574gat | n1573gat;
assign n2992gat = n1723gat | n1647gat | n1646gat;
assign n2986gat = n1650gat | n1649gat | n1563gat;
assign n2991gat = n1654gat | n1653gat | n1644gat;
assign II3148 = n1839gat | n1884gat | n1784gat;
assign II3149 = n1786gat | n1787gat | II3148;
assign II3178 = n1838gat | n1785gat | n1788gat;
assign II3179 = n1839gat | n1784gat | II3178;
assign n2981gat = n1413gat | n1408gat | n1407gat;
assign n3000gat = n2000gat | n1999gat;
assign n3004gat = n2258gat | n2257gat | n2255gat;
assign n3003gat = n2256gat | n2251gat;
assign n3001gat = n2132gat | n2130gat;
assign n3006gat = n2253gat | n2252gat;
assign n3007gat = n2250gat | n2249gat;
assign n2990gat = n1710gat | n1630gat;
assign n2994gat = n1954gat | n1888gat;
assign n2993gat = n1894gat | n1847gat | n1846gat;
assign n2998gat = n2055gat | n1967gat;
assign n2996gat = n1960gat | n1959gat | n1957gat;
assign n3008gat = n2332gat | n2259gat;
assign n3005gat = n2211gat | n2210gat;
assign n2997gat = n2053gat | n2052gat | n1964gat;
assign n3009gat = n2350gat | n2282gat;
assign n3002gat = n2213gat | n2150gat | n2149gat;
assign n2995gat = n1962gat | n1955gat;
assign n2999gat = n1972gat | n1971gat;
assign n3011gat = n2333gat | n2331gat;
assign n3015gat = n2566gat | n2565gat;
assign n2874gat = n141gat | n38gat | n37gat;
assign n2917gat = n1074gat | n872gat;
assign n2878gat = n234gat | n137gat;
assign n2892gat = n378gat | n377gat;
assign n2885gat = n250gat | n249gat | n248gat;
assign n2900gat = n869gat | n453gat | n448gat;
assign n2883gat = n251gat | n244gat;
assign n2929gat = n974gat | n973gat | n870gat;
assign n2884gat = n246gat | n245gat;
assign n2902gat = n460gat | n459gat;
assign n2925gat = n975gat | n972gat | n969gat;
assign n2879gat = n145gat | n143gat;
assign n2916gat = n971gat | n970gat | n968gat;
assign n2875gat = n142gat | n40gat | n39gat;
assign n2899gat = n772gat | n451gat | n446gat;
assign n2877gat = n139gat | n136gat;
assign n2893gat = n391gat | n390gat;
assign n2926gat = n1083gat | n1077gat;
assign n2882gat = n242gat | n240gat;
assign n2924gat = n871gat | n797gat;
assign n2881gat = n324gat | n238gat | n237gat;
assign n2923gat = n1082gat | n796gat;
assign n2710gat = n69gat | n1885gat;
assign n2704gat = n11gat | n1889gat;
assign n2684gat = n1599gat | n2051gat;
assign n2830gat = n2444gat | n1754gat;
assign II3999 = n2167gat | n2031gat | n2174gat;
assign II4000 = n2108gat | n2093gat | n2035gat | II3999;
assign n2695gat = n1586gat | n1791gat;
assign n2703gat = n1755gat | n1518gat;
assign n2744gat = n2159gat | n2478gat;
assign n2800gat = n2158gat | n2186gat;
assign II4023 = n2443gat | n2290gat | n2214gat;
assign II4024 = n2353gat | n2284gat | II4023;
assign n2980gat = n1470gat | n1400gat | n1399gat | n1398gat;
assign II4144 = n1633gat | n1838gat | n1786gat;
assign II4145 = n1788gat | n1784gat | II4144;
assign n2984gat = n1467gat | n1466gat;
assign n2985gat = n1686gat | n1533gat | n1532gat | n1531gat;
assign II4216 = n1427gat | n1595gat | n1677gat;
assign II4217 = n1392gat | n2989gat | II4216;
assign n2931gat = n1100gat | n994gat | n989gat | n880gat;
assign n2943gat = n1012gat | n905gat;
assign n2941gat = n1003gat | n902gat;
assign n2946gat = n1099gat | n998gat | n995gat | n980gat;
assign n2960gat = n1175gat | n1174gat;
assign n2950gat = n1001gat | n999gat;
assign n2969gat = n1323gat | n1264gat;
assign n2933gat = n981gat | n890gat | n889gat | n886gat;
assign n2935gat = n892gat | n891gat;
assign n2942gat = n904gat | n903gat;
assign n2940gat = n1152gat | n1092gat | n997gat | n993gat;
assign n2937gat = n900gat | n895gat;
assign n2947gat = n1094gat | n1093gat | n988gat | n984gat;
assign n2965gat = n1267gat | n1257gat;
assign n2956gat = n1178gat | n1116gat;
assign n2961gat = n1375gat | n1324gat;
assign n2939gat = n1091gat | n1088gat | n992gat | n987gat;
assign n2938gat = n899gat | n896gat;
assign n2967gat = n1262gat | n1260gat;
assign n2932gat = n1098gat | n1090gat | n986gat | n885gat;
assign n2936gat = n901gat | n893gat;
assign n2948gat = n1097gat | n1089gat | n1087gat | n991gat;
assign n2968gat = n1326gat | n1261gat;
assign n2955gat = n1177gat | n1115gat;
assign n2944gat = n977gat | n976gat;
assign n2945gat = n1096gat | n1095gat | n990gat | n979gat;
assign n2962gat = n1176gat | n1173gat;
assign n2951gat = n1004gat | n1000gat;
assign n2764gat = n1029gat | n2237gat;
assign n2762gat = n1028gat | n1782gat;
assign n2761gat = n1031gat | n2325gat;
assign n2757gat = n1030gat | n2245gat;
assign n2756gat = n1011gat | n2244gat;
assign n2750gat = n1181gat | n2243gat;
assign n2749gat = n1010gat | n2246gat;
assign n2742gat = n1005gat | n2384gat;
assign n2741gat = n1182gat | n2385gat;
assign n2694gat = n1381gat | n1384gat;
assign n2693gat = n1451gat | n1453gat;
assign n2702gat = n925gat | n1452gat;
assign n2701gat = n921gat | n1890gat;
assign n2709gat = n739gat | n1841gat;
assign n2708gat = n848gat | n2047gat;
assign n2799gat = n849gat | n2050gat;
assign n2798gat = n1032gat | n2054gat;
assign n2812gat = n73gat | n70gat | n1840gat;
assign n2822gat = n77gat | n13gat | n1842gat;
assign n421gat = ~(n2715gat | n2723gat);
assign n648gat = ~(n373gat | n2669gat);
assign n442gat = ~(n2844gat | n856gat);
assign n1499gat = ~(n396gat | n401gat);
assign n1616gat = ~(n918gat | n396gat);
assign n1614gat = ~(n396gat | n845gat);
assign n1641gat = ~(n1645gat | n1553gat | n1559gat);
assign n1642gat = ~(n1559gat | n1616gat | n1645gat);
assign n1556gat = ~(n1614gat | n1645gat | n1616gat);
assign n1557gat = ~(n1553gat | n1645gat | n1614gat);
assign n1639gat = ~(n1499gat | n1559gat | n1553gat);
assign n1605gat = ~(n1614gat | n1616gat | n1499gat | n396gat);
assign n1555gat = ~(n1616gat | n1559gat | n1499gat);
assign n1558gat = ~(n1614gat | n1553gat | n1499gat);
assign n1256gat = ~(n392gat | n702gat);
assign n1117gat = ~(n720gat | n725gat);
assign n1618gat = ~(n1319gat | n1447gat);
assign n1114gat = ~(n725gat | n721gat);
assign n1621gat = ~(n1319gat | n1380gat);
assign n1318gat = ~(n392gat | n701gat);
assign n1619gat = ~(n1447gat | n1446gat);
assign n1622gat = ~(n1380gat | n1446gat);
assign n1214gat = ~(n1218gat | n1219gat | n1220gat);
assign n1215gat = ~(n1218gat | n1221gat | n1222gat);
assign n1216gat = ~(n1223gat | n1219gat | n1222gat);
assign n1217gat = ~(n1223gat | n1221gat | n1220gat);
assign n745gat = ~(n2716gat | n2867gat);
assign n638gat = ~(n2715gat | n2868gat);
assign n423gat = ~(n2724gat | n2726gat);
assign n362gat = ~(n2723gat | n2727gat);
assign n749gat = ~(n753gat | n754gat | n755gat);
assign n750gat = ~(n753gat | n756gat | n757gat);
assign n751gat = ~(n758gat | n754gat | n757gat);
assign n752gat = ~(n758gat | n756gat | n755gat);
assign n259gat = ~(n263gat | n264gat | n265gat);
assign n260gat = ~(n263gat | n266gat | n267gat);
assign n261gat = ~(n268gat | n264gat | n267gat);
assign n262gat = ~(n268gat | n266gat | n265gat);
assign n1014gat = ~(n1018gat | n1019gat | n1020gat);
assign n1015gat = ~(n1018gat | n1021gat | n1022gat);
assign n1016gat = ~(n1023gat | n1019gat | n1022gat);
assign n1017gat = ~(n1023gat | n1021gat | n1020gat);
assign n476gat = ~(n480gat | n481gat | n482gat);
assign n477gat = ~(n480gat | n483gat | n484gat);
assign n478gat = ~(n485gat | n481gat | n484gat);
assign n479gat = ~(n485gat | n483gat | n482gat);
assign n44gat = ~(n48gat | n49gat | n50gat);
assign n45gat = ~(n48gat | n51gat | n52gat);
assign n46gat = ~(n53gat | n49gat | n52gat);
assign n47gat = ~(n53gat | n51gat | n50gat);
assign n1376gat = ~(n724gat | n720gat);
assign n1617gat = ~(n1319gat | n1448gat);
assign n1377gat = ~(n724gat | n721gat);
assign n1624gat = ~(n1319gat | n1379gat);
assign n1113gat = ~(n393gat | n701gat);
assign n1501gat = ~(n1448gat | n1500gat);
assign n1623gat = ~(n1379gat | n1446gat);
assign n1620gat = ~(n1448gat | n1446gat);
assign n1827gat = ~(n2729gat | n2317gat);
assign n1817gat = ~(n1819gat | n1823gat);
assign n1935gat = ~(n1816gat | n1828gat);
assign n529gat = ~(n2724gat | n2715gat);
assign n361gat = ~(n2859gat | n2726gat);
assign n168gat = ~(n172gat | n173gat | n174gat);
assign n169gat = ~(n172gat | n175gat | n176gat);
assign n170gat = ~(n177gat | n173gat | n176gat);
assign n171gat = ~(n177gat | n175gat | n174gat);
assign n907gat = ~(n911gat | n912gat | n913gat);
assign n908gat = ~(n911gat | n914gat | n915gat);
assign n909gat = ~(n916gat | n912gat | n915gat);
assign n910gat = ~(n916gat | n914gat | n913gat);
assign n344gat = ~(n348gat | n349gat | n350gat);
assign n345gat = ~(n348gat | n351gat | n352gat);
assign n346gat = ~(n353gat | n349gat | n352gat);
assign n347gat = ~(n353gat | n351gat | n350gat);
assign n56gat = ~(n60gat | n61gat | n62gat);
assign n57gat = ~(n60gat | n63gat | n64gat);
assign n58gat = ~(n65gat | n61gat | n64gat);
assign n59gat = ~(n65gat | n63gat | n62gat);
assign n768gat = ~(n373gat | n2731gat);
assign n655gat = ~(n856gat | n2718gat);
assign n963gat = ~(n856gat | n2838gat);
assign n868gat = ~(n2775gat | n373gat);
assign n962gat = ~(n856gat | n2711gat);
assign n959gat = ~(n373gat | n2734gat);
assign n945gat = ~(n949gat | n950gat | n951gat);
assign n946gat = ~(n949gat | n952gat | n953gat);
assign n947gat = ~(n954gat | n950gat | n953gat);
assign n948gat = ~(n954gat | n952gat | n951gat);
assign n647gat = ~(n2792gat | n373gat);
assign n441gat = ~(n856gat | n2846gat);
assign n967gat = ~(n373gat | n2672gat);
assign n792gat = ~(n2852gat | n856gat);
assign n1229gat = ~(n1233gat | n1234gat | n1235gat);
assign n1230gat = ~(n1233gat | n1236gat | n1237gat);
assign n1231gat = ~(n1238gat | n1234gat | n1237gat);
assign n1232gat = ~(n1238gat | n1236gat | n1235gat);
assign n443gat = ~(n2778gat | n373gat);
assign n439gat = ~(n856gat | n2836gat);
assign n966gat = ~(n2789gat | n373gat);
assign n790gat = ~(n856gat | n2840gat);
assign n444gat = ~(n373gat | n2781gat);
assign n440gat = ~(n856gat | n2842gat);
assign n1051gat = ~(n1055gat | n1056gat | n1057gat);
assign n1052gat = ~(n1055gat | n1058gat | n1059gat);
assign n1053gat = ~(n1060gat | n1056gat | n1059gat);
assign n1054gat = ~(n1060gat | n1058gat | n1057gat);
assign n934gat = ~(n938gat | n939gat | n940gat);
assign n935gat = ~(n938gat | n941gat | n942gat);
assign n936gat = ~(n943gat | n939gat | n942gat);
assign n937gat = ~(n943gat | n941gat | n940gat);
assign n746gat = ~(n2716gat | n2723gat);
assign n360gat = ~(n2859gat | n2727gat);
assign n710gat = ~(n714gat | n715gat | n716gat);
assign n711gat = ~(n714gat | n717gat | n718gat);
assign n712gat = ~(n719gat | n715gat | n718gat);
assign n713gat = ~(n719gat | n717gat | n716gat);
assign n729gat = ~(n733gat | n734gat | n735gat);
assign n730gat = ~(n733gat | n736gat | n737gat);
assign n731gat = ~(n738gat | n734gat | n737gat);
assign n732gat = ~(n738gat | n736gat | n735gat);
assign n494gat = ~(n498gat | n499gat | n500gat);
assign n495gat = ~(n498gat | n501gat | n502gat);
assign n496gat = ~(n503gat | n499gat | n502gat);
assign n497gat = ~(n503gat | n501gat | n500gat);
assign n505gat = ~(n509gat | n510gat | n511gat);
assign n506gat = ~(n509gat | n512gat | n513gat);
assign n507gat = ~(n514gat | n510gat | n513gat);
assign n508gat = ~(n514gat | n512gat | n511gat);
assign n564gat = ~(n3029gat | n2863gat | n2855gat | n374gat);
assign n86gat = ~(n743gat | n294gat | n17gat);
assign n78gat = ~(n2784gat | n79gat);
assign n767gat = ~(n219gat | n2731gat);
assign n286gat = ~(n289gat | n2723gat);
assign n287gat = ~(n289gat | n2715gat);
assign n288gat = ~(n289gat | n2726gat);
assign n181gat = ~(n286gat | n179gat | n188gat);
assign n182gat = ~(n72gat | n2720gat);
assign n653gat = ~(n2718gat | n111gat);
assign n867gat = ~(n219gat | n2775gat);
assign n771gat = ~(n2838gat | n111gat);
assign n964gat = ~(n111gat | n2711gat);
assign n961gat = ~(n219gat | n2734gat);
assign n804gat = ~(n808gat | n809gat | n810gat);
assign n805gat = ~(n808gat | n811gat | n812gat);
assign n806gat = ~(n813gat | n809gat | n812gat);
assign n807gat = ~(n813gat | n811gat | n810gat);
assign n587gat = ~(n591gat | n592gat | n593gat);
assign n588gat = ~(n591gat | n594gat | n595gat);
assign n589gat = ~(n596gat | n592gat | n595gat);
assign n590gat = ~(n596gat | n594gat | n593gat);
assign n447gat = ~(n2836gat | n111gat);
assign n445gat = ~(n2778gat | n219gat);
assign n687gat = ~(n691gat | n692gat | n693gat);
assign n688gat = ~(n691gat | n694gat | n695gat);
assign n689gat = ~(n696gat | n692gat | n695gat);
assign n690gat = ~(n696gat | n694gat | n693gat);
assign n568gat = ~(n572gat | n573gat | n574gat);
assign n569gat = ~(n572gat | n575gat | n576gat);
assign n570gat = ~(n577gat | n573gat | n576gat);
assign n571gat = ~(n577gat | n575gat | n574gat);
assign n187gat = ~(n189gat | n287gat | n188gat);
assign n197gat = ~(n194gat | n297gat);
assign n15gat = ~(n637gat | n17gat | n293gat);
assign n22gat = ~(n92gat | n21gat);
assign n93gat = ~(n197gat | n22gat);
assign n769gat = ~(n93gat | n2731gat);
assign n2534gat = ~(n2624gat | n2489gat | n2621gat);
assign n2430gat = ~(n2533gat | n2486gat | n2429gat);
assign n1606gat = ~(n3020gat | n270gat);
assign n2239gat = ~(n2850gat | n3019gat);
assign n1934gat = ~(n2470gat | n1935gat | n2239gat);
assign n1610gat = ~(n1698gat | n1543gat);
assign n1692gat = ~(n1879gat | n1762gat);
assign n2433gat = ~(n2432gat | n2154gat);
assign n2531gat = ~(n2488gat | n2625gat | n2621gat);
assign n2480gat = ~(n2530gat | n2482gat | n2486gat);
assign n2427gat = ~(n2426gat | n2153gat);
assign n2428gat = ~(n2433gat | n2427gat);
assign n1778gat = ~(n3026gat | n1779gat);
assign n1609gat = ~(n1503gat | n3025gat);
assign n1702gat = ~(n3024gat | n1615gat);
assign n1700gat = ~(n1701gat | n3023gat);
assign n1604gat = ~(n1778gat | n1609gat | n1702gat | n1700gat);
assign n1076gat = ~(n93gat | n2775gat);
assign n766gat = ~(n93gat | n2734gat);
assign n1185gat = ~(n1189gat | n1190gat | n1191gat);
assign n1186gat = ~(n1189gat | n1192gat | n1193gat);
assign n1187gat = ~(n1194gat | n1190gat | n1193gat);
assign n1188gat = ~(n1194gat | n1192gat | n1191gat);
assign n645gat = ~(n2792gat | n93gat);
assign n646gat = ~(n93gat | n2669gat);
assign n1383gat = ~(n1280gat | n1225gat);
assign n1327gat = ~(n1281gat | n1224gat);
assign n651gat = ~(n93gat | n2778gat);
assign n652gat = ~(n2789gat | n93gat);
assign n765gat = ~(n2781gat | n93gat);
assign n1202gat = ~(n1206gat | n1207gat | n1208gat);
assign n1203gat = ~(n1206gat | n1209gat | n1210gat);
assign n1204gat = ~(n1211gat | n1207gat | n1210gat);
assign n1205gat = ~(n1211gat | n1209gat | n1208gat);
assign n1270gat = ~(n1274gat | n1275gat | n1276gat);
assign n1271gat = ~(n1274gat | n1277gat | n1278gat);
assign n1272gat = ~(n1279gat | n1275gat | n1278gat);
assign n1273gat = ~(n1279gat | n1277gat | n1276gat);
assign n763gat = ~(n2672gat | n93gat);
assign n1287gat = ~(n1284gat | n1195gat);
assign n1285gat = ~(n1196gat | n1269gat);
assign n853gat = ~(n740gat | n2148gat);
assign n793gat = ~(n2852gat | n851gat);
assign n854gat = ~(n2148gat | n374gat);
assign n556gat = ~(n2672gat | n852gat);
assign n795gat = ~(n2731gat | n852gat);
assign n656gat = ~(n851gat | n2718gat);
assign n794gat = ~(n852gat | n2775gat);
assign n773gat = ~(n851gat | n2838gat);
assign n965gat = ~(n2711gat | n851gat);
assign n960gat = ~(n2734gat | n852gat);
assign n780gat = ~(n784gat | n785gat | n786gat);
assign n781gat = ~(n784gat | n787gat | n788gat);
assign n782gat = ~(n789gat | n785gat | n788gat);
assign n783gat = ~(n789gat | n787gat | n786gat);
assign n555gat = ~(n852gat | n2792gat);
assign n450gat = ~(n851gat | n2846gat);
assign n654gat = ~(n851gat | n2844gat);
assign n557gat = ~(n2669gat | n852gat);
assign n874gat = ~(n559gat | n365gat);
assign n132gat = ~(n560gat | n364gat);
assign n649gat = ~(n2778gat | n852gat);
assign n449gat = ~(n2836gat | n851gat);
assign n791gat = ~(n851gat | n2840gat);
assign n650gat = ~(n852gat | n2789gat);
assign n774gat = ~(n2842gat | n851gat);
assign n764gat = ~(n852gat | n2781gat);
assign n222gat = ~(n226gat | n227gat | n228gat);
assign n223gat = ~(n226gat | n229gat | n230gat);
assign n224gat = ~(n231gat | n227gat | n230gat);
assign n225gat = ~(n231gat | n229gat | n228gat);
assign n121gat = ~(n125gat | n126gat | n127gat);
assign n122gat = ~(n125gat | n128gat | n129gat);
assign n123gat = ~(n130gat | n126gat | n129gat);
assign n124gat = ~(n130gat | n128gat | n127gat);
assign n2460gat = ~(n666gat | n120gat);
assign n2423gat = ~(n665gat | n1601gat);
assign n2594gat = ~(n3017gat | n2520gat | n2597gat);
assign n2569gat = ~(n2573gat | n2574gat | n2575gat);
assign n2570gat = ~(n2573gat | n2576gat | n2577gat);
assign n2571gat = ~(n2578gat | n2574gat | n2577gat);
assign n2572gat = ~(n2578gat | n2576gat | n2575gat);
assign n2410gat = ~(n2414gat | n2415gat | n2416gat);
assign n2411gat = ~(n2414gat | n2417gat | n2418gat);
assign n2412gat = ~(n2419gat | n2415gat | n2418gat);
assign n2413gat = ~(n2419gat | n2417gat | n2416gat);
assign n2583gat = ~(n2582gat | n2585gat);
assign n2580gat = ~(n2582gat | n2583gat);
assign n2581gat = ~(n2583gat | n2585gat);
assign n2567gat = ~(n2493gat | n2388gat);
assign n2499gat = ~(n2389gat | n2494gat);
assign n299gat = ~(n2268gat | n2338gat);
assign n207gat = ~(n2337gat | n2269gat);
assign n2650gat = ~(n2649gat | n2652gat);
assign n2647gat = ~(n2649gat | n2650gat);
assign n2648gat = ~(n2650gat | n2652gat);
assign n2602gat = ~(n2606gat | n2607gat | n2608gat);
assign n2603gat = ~(n2606gat | n2609gat | n2610gat);
assign n2604gat = ~(n2611gat | n2607gat | n2610gat);
assign n2605gat = ~(n2611gat | n2609gat | n2608gat);
assign n2546gat = ~(n2550gat | n2551gat | n2552gat);
assign n2547gat = ~(n2550gat | n2553gat | n2554gat);
assign n2548gat = ~(n2555gat | n2551gat | n2554gat);
assign n2549gat = ~(n2555gat | n2553gat | n2552gat);
assign n2617gat = ~(n2616gat | n2619gat);
assign n2614gat = ~(n2616gat | n2617gat);
assign n2615gat = ~(n2617gat | n2619gat);
assign n2655gat = ~(n2508gat | n2656gat | n2500gat | n2504gat);
assign n2293gat = ~(n2353gat | n2284gat | n2443gat);
assign n2219gat = ~(n2354gat | n2214gat);
assign n1529gat = ~(n1528gat | n1523gat);
assign n1704gat = ~(n3027gat | n1706gat);
assign n2461gat = ~(n120gat | n2666gat);
assign n2421gat = ~(n1601gat | n1704gat);
assign n1598gat = ~(n1592gat | n2422gat);
assign n2218gat = ~(n2214gat | n2290gat);
assign n2358gat = ~(n2285gat | n2356gat | n2355gat);
assign n1415gat = ~(n2081gat | n2359gat);
assign n1153gat = ~(n1414gat | n566gat);
assign n2292gat = ~(n2443gat | n2284gat | n2285gat);
assign n1416gat = ~(n2081gat | n1480gat);
assign n1151gat = ~(n1301gat | n1150gat);
assign n2306gat = ~(n2356gat | n2284gat | n2285gat);
assign n1481gat = ~(n2081gat | n2011gat);
assign n982gat = ~(n873gat | n1478gat);
assign n2357gat = ~(n2285gat | n2355gat | n2443gat);
assign n1347gat = ~(n2081gat | n1410gat);
assign n877gat = ~(n875gat | n876gat);
assign n1484gat = ~(n2081gat | n1528gat);
assign n1159gat = ~(n1160gat | n1084gat);
assign n2363gat = ~(n2353gat | n2356gat | n2355gat);
assign n1483gat = ~(n2081gat | n1482gat);
assign n1158gat = ~(n983gat | n1157gat);
assign n2364gat = ~(n2353gat | n2284gat | n2356gat);
assign n1308gat = ~(n2081gat | n1530gat);
assign n1156gat = ~(n985gat | n1307gat);
assign n2291gat = ~(n2353gat | n2355gat | n2443gat);
assign n1349gat = ~(n1479gat | n2081gat);
assign n1155gat = ~(n1085gat | n1348gat);
assign n1154gat = ~(n1598gat | n2930gat | n2957gat);
assign n1703gat = ~(n1705gat | n3028gat);
assign n1608gat = ~(n1704gat | n1703gat);
assign n1411gat = ~(n1154gat | n1608gat);
assign n2223gat = ~(n2354gat | n2217gat);
assign n1438gat = ~(n1591gat | n1480gat);
assign n1625gat = ~(n3021gat | n1628gat);
assign n1626gat = ~(n1627gat | n3022gat);
assign n1831gat = ~(n1832gat | n1765gat | n1878gat);
assign n1443gat = ~(n1442gat | n706gat);
assign n1325gat = ~(n1444gat | n164gat);
assign n1441gat = ~(n1437gat | n1378gat);
assign n1321gat = ~(n1442gat | n837gat);
assign n1320gat = ~(n1444gat | n278gat);
assign n1486gat = ~(n1482gat | n1591gat);
assign n1440gat = ~(n1322gat | n1439gat);
assign n1426gat = ~(n2011gat | n1591gat);
assign n1368gat = ~(n1442gat | n613gat);
assign n1258gat = ~(n274gat | n1444gat);
assign n1371gat = ~(n1370gat | n1369gat);
assign n1365gat = ~(n1479gat | n1591gat);
assign n1373gat = ~(n833gat | n1442gat);
assign n1372gat = ~(n282gat | n1444gat);
assign n1367gat = ~(n1366gat | n1374gat);
assign n2220gat = ~(n2290gat | n2217gat);
assign n1423gat = ~(n2162gat | n1530gat);
assign n1498gat = ~(n1609gat | n1427gat);
assign n1504gat = ~(n1450gat | n1498gat);
assign n1607gat = ~(n2082gat | n1609gat);
assign n1494gat = ~(n1528gat | n2162gat);
assign n1502gat = ~(n1607gat | n1449gat);
assign n1250gat = ~(n1603gat | n815gat);
assign n1103gat = ~(n956gat | n1590gat);
assign n1417gat = ~(n2162gat | n1480gat);
assign n1352gat = ~(n1248gat | n1418gat);
assign n1304gat = ~(n1590gat | n1067gat);
assign n1249gat = ~(n679gat | n1603gat);
assign n1419gat = ~(n2162gat | n1479gat);
assign n1351gat = ~(n1306gat | n1353gat);
assign n1246gat = ~(n864gat | n1590gat);
assign n1161gat = ~(n583gat | n1603gat);
assign n1422gat = ~(n2011gat | n2162gat);
assign n1303gat = ~(n1247gat | n1355gat);
assign n1291gat = ~(n1603gat | n579gat);
assign n1245gat = ~(n1590gat | n860gat);
assign n1485gat = ~(n1482gat | n2162gat);
assign n1302gat = ~(n1300gat | n1487gat);
assign n1163gat = ~(n882gat | n1603gat);
assign n1102gat = ~(n1297gat | n1590gat);
assign n1354gat = ~(n1591gat | n1530gat);
assign n1360gat = ~(n1164gat | n1356gat);
assign n1435gat = ~(n1591gat | n1528gat);
assign n1101gat = ~(n1590gat | n1293gat);
assign n996gat = ~(n1603gat | n823gat);
assign n1359gat = ~(n1436gat | n1106gat);
assign n1421gat = ~(n2162gat | n2359gat);
assign n1104gat = ~(n1079gat | n1590gat);
assign n887gat = ~(n1603gat | n683gat);
assign n1358gat = ~(n1425gat | n1105gat);
assign n1420gat = ~(n1410gat | n2162gat);
assign n1305gat = ~(n1147gat | n1590gat);
assign n1162gat = ~(n698gat | n1603gat);
assign n1357gat = ~(n1424gat | n1309gat);
assign n1428gat = ~(n2978gat | n2982gat | n2973gat | n2977gat);
assign n1794gat = ~(n1673gat | n1719gat);
assign n1796gat = ~(n1858gat | n1635gat);
assign n1792gat = ~(n1794gat | n1796gat);
assign n1865gat = ~(n1989gat | n1918gat | n1986gat);
assign n1861gat = ~(n1866gat | n2216gat | n1988gat);
assign n1793gat = ~(n1792gat | n1735gat);
assign n1406gat = ~(n1428gat | n1387gat);
assign n1780gat = ~(n1777gat | n1625gat | n1626gat);
assign n2016gat = ~(n2019gat | n1878gat);
assign n2664gat = ~(n2850gat | n3018gat);
assign n1666gat = ~(n1986gat | n2212gat | n1991gat);
assign n1578gat = ~(n2152gat | n2351gat | n1665gat);
assign n1516gat = ~(n1551gat | n1517gat);
assign n1864gat = ~(n1858gat | n1495gat | n2090gat);
assign n1565gat = ~(n1735gat | n1552gat);
assign n1921gat = ~(n1738gat | n1673gat);
assign n1798gat = ~(n1739gat | n1673gat);
assign n1920gat = ~(n1864gat | n1921gat | n1798gat);
assign n1926gat = ~(n1925gat | n1635gat);
assign n1916gat = ~(n1917gat | n1859gat);
assign n1994gat = ~(n1719gat | n1922gat);
assign n1924gat = ~(n1743gat | n1923gat);
assign n2078gat = ~(n1926gat | n1916gat | n1994gat | n1924gat);
assign n1690gat = ~(n1700gat | n1702gat);
assign n1660gat = ~(n1918gat | n1986gat | n2212gat);
assign n1576gat = ~(n2351gat | n1988gat | n1661gat);
assign n1733gat = ~(n1673gat | n1572gat);
assign n1582gat = ~(n2283gat | n1991gat | n2212gat);
assign n1577gat = ~(n1520gat | n2351gat | n1988gat);
assign n1581gat = ~(n1858gat | n1580gat);
assign n2129gat = ~(n2189gat | n2134gat | n2261gat);
assign n2079gat = ~(n2078gat | n2178gat | n1990gat | n2128gat);
assign n1695gat = ~(n1609gat | n1778gat | n1704gat | n1703gat);
assign n2073gat = ~(n2078gat | n1990gat | n2181gat);
assign n1696gat = ~(n1707gat | n1698gat);
assign n1758gat = ~(n1311gat | n1773gat);
assign n1574gat = ~(n1719gat | n1673gat | n1444gat);
assign n1573gat = ~(n1444gat | n1858gat | n1635gat);
assign n1521gat = ~(n2283gat | n1991gat);
assign n1737gat = ~(n2212gat | n2152gat);
assign n1732gat = ~(n1515gat | n1736gat | n1658gat);
assign n1723gat = ~(n1659gat | n1722gat | n1724gat);
assign n1663gat = ~(n1986gat | n1918gat);
assign n1655gat = ~(n1736gat | n1662gat | n1658gat);
assign n1647gat = ~(n1656gat | n1659gat | n1554gat);
assign n1667gat = ~(n1991gat | n1986gat);
assign n1570gat = ~(n1736gat | n1658gat | n1670gat);
assign n1646gat = ~(n1569gat | n1659gat | n1566gat);
assign n1575gat = ~(n1918gat | n2283gat);
assign n1728gat = ~(n1568gat | n1736gat | n1658gat);
assign n1650gat = ~(n1727gat | n1659gat | n1640gat);
assign n1801gat = ~(n2152gat | n1989gat);
assign n1731gat = ~(n1658gat | n1515gat | n1797gat);
assign n1649gat = ~(n1560gat | n1659gat | n1730gat);
assign n1571gat = ~(n1670gat | n1658gat | n1797gat);
assign n1563gat = ~(n1561gat | n1562gat | n1659gat);
assign n1734gat = ~(n1988gat | n2212gat);
assign n1669gat = ~(n1668gat | n1742gat | n1670gat);
assign n1654gat = ~(n1671gat | n1659gat);
assign n1657gat = ~(n1662gat | n1797gat | n1658gat);
assign n1653gat = ~(n1651gat | n1652gat | n1659gat);
assign n1729gat = ~(n1658gat | n1797gat | n1568gat);
assign n1644gat = ~(n1643gat | n1648gat | n1659gat);
assign n1726gat = ~(n2992gat | n2986gat | n2991gat);
assign n1929gat = ~(n1758gat | n1790gat);
assign n2009gat = ~(n2016gat | n2664gat | n2004gat);
assign n1413gat = ~(n1869gat | n672gat | n2591gat);
assign n1636gat = ~(n1584gat | n1718gat);
assign n1401gat = ~(n1584gat | n1590gat);
assign n1408gat = ~(n1507gat | n1396gat | n1393gat);
assign n1476gat = ~(n1858gat | n1590gat);
assign n1407gat = ~(n1393gat | n1409gat | n1677gat);
assign n1412gat = ~(n1411gat | n1406gat | n2981gat);
assign n2663gat = ~(n2586gat | n2660gat | n2307gat);
assign n2662gat = ~(n2660gat | n2586gat);
assign n2238gat = ~(n2448gat | n2444gat);
assign n87gat = ~(n743gat | n17gat | n293gat);
assign n200gat = ~(n199gat | n92gat);
assign n184gat = ~(n189gat | n188gat | n179gat);
assign n196gat = ~(n297gat | n195gat);
assign n204gat = ~(n200gat | n196gat);
assign n2163gat = ~(n1790gat | n1310gat | n2664gat | n2168gat);
assign n2258gat = ~(n2260gat | n2189gat);
assign n2255gat = ~(n2261gat | n2188gat);
assign n2015gat = ~(n2039gat | n1774gat | n1315gat);
assign n2017gat = ~(n1790gat | n2016gat);
assign n2018gat = ~(n2016gat | n2097gat);
assign n2014gat = ~(n2035gat | n2093gat | n2018gat | n2664gat);
assign n2194gat = ~(n2187gat | n1855gat);
assign n2192gat = ~(n2184gat | n1855gat);
assign n2185gat = ~(n2261gat | n2189gat);
assign n2132gat = ~(n2133gat | n2131gat);
assign n2130gat = ~(n2134gat | n2185gat);
assign n2057gat = ~(n2049gat | n1855gat);
assign n2250gat = ~(n2248gat | n2264gat);
assign n2249gat = ~(n2265gat | n3006gat);
assign n2329gat = ~(n1855gat | n3007gat);
assign n1958gat = ~(n1963gat | n1886gat);
assign n1895gat = ~(n1845gat | n1891gat | n1968gat);
assign n1710gat = ~(n1709gat | n1629gat);
assign n1630gat = ~(n1895gat | n1631gat);
assign n2195gat = ~(n2200gat | n1855gat);
assign n2556gat = ~(n1711gat | n2437gat);
assign n2539gat = ~(n2048gat | n2437gat);
assign n1894gat = ~(n1968gat | n1891gat | n1969gat);
assign n1847gat = ~(n1958gat | n1845gat);
assign n1846gat = ~(n1845gat | n1893gat);
assign n2436gat = ~(n2437gat | n1892gat);
assign n2055gat = ~(n1891gat | n1958gat);
assign n1967gat = ~(n1893gat | n1968gat);
assign n2387gat = ~(n2056gat | n2437gat);
assign n1959gat = ~(n1956gat | n1963gat);
assign n1957gat = ~(n1886gat | n1887gat);
assign n2330gat = ~(n2437gat | n1961gat);
assign n2147gat = ~(n2988gat | n1855gat);
assign n2498gat = ~(n2199gat | n2328gat);
assign n2193gat = ~(n2393gat | n2439gat);
assign n2211gat = ~(n2193gat | n2402gat);
assign n2210gat = ~(n2401gat | n2151gat);
assign n2396gat = ~(n2199gat | n2209gat);
assign n2053gat = ~(n2393gat | n2438gat);
assign n1964gat = ~(n2392gat | n2439gat);
assign n2198gat = ~(n2199gat | n2058gat);
assign n2215gat = ~(n2346gat | n2151gat | n2402gat);
assign n2350gat = ~(n2405gat | n2349gat);
assign n2282gat = ~(n2406gat | n2215gat);
assign n2197gat = ~(n2199gat | n2281gat);
assign n2213gat = ~(n2402gat | n2151gat | n2345gat);
assign n2150gat = ~(n2401gat | n2346gat);
assign n2149gat = ~(n2193gat | n2346gat);
assign n2196gat = ~(n2199gat | n2146gat);
assign n1882gat = ~(n2124gat | n2115gat | n2239gat);
assign n1962gat = ~(n1963gat | n1893gat);
assign n1896gat = ~(n2995gat | n1895gat);
assign n1972gat = ~(n1974gat | n1970gat);
assign n1971gat = ~(n1896gat | n1973gat);
assign n2559gat = ~(n2999gat | n2437gat);
assign n2331gat = ~(n2393gat | n2401gat);
assign n2352gat = ~(n3011gat | n2215gat);
assign n2566gat = ~(n2643gat | n2564gat);
assign n2565gat = ~(n2352gat | n2642gat);
assign n2637gat = ~(n3015gat | n2199gat);
assign n84gat = ~(n296gat | n17gat | n294gat);
assign n89gat = ~(n88gat | n2784gat);
assign n110gat = ~(n182gat | n89gat);
assign n1074gat = ~(n2775gat | n110gat);
assign n141gat = ~(n155gat | n253gat | n150gat);
assign n38gat = ~(n151gat | n233gat);
assign n37gat = ~(n151gat | n154gat);
assign n872gat = ~(n375gat | n800gat);
assign n234gat = ~(n155gat | n233gat);
assign n137gat = ~(n154gat | n253gat);
assign n378gat = ~(n375gat | n235gat);
assign n377gat = ~(n110gat | n2778gat);
assign n869gat = ~(n219gat | n2792gat);
assign n212gat = ~(n182gat | n78gat);
assign n250gat = ~(n329gat | n387gat | n334gat);
assign n249gat = ~(n386gat | n330gat);
assign n248gat = ~(n330gat | n1490gat);
assign n453gat = ~(n372gat | n452gat);
assign n448gat = ~(n111gat | n2846gat);
assign n974gat = ~(n2844gat | n111gat);
assign n251gat = ~(n1490gat | n387gat);
assign n244gat = ~(n334gat | n386gat);
assign n973gat = ~(n372gat | n333gat);
assign n870gat = ~(n2669gat | n219gat);
assign n975gat = ~(n111gat | n2852gat);
assign n246gat = ~(n330gat | n325gat | n334gat);
assign n245gat = ~(n386gat | n334gat);
assign n460gat = ~(n462gat | n2884gat);
assign n459gat = ~(n457gat | n461gat);
assign n972gat = ~(n372gat | n458gat);
assign n969gat = ~(n219gat | n2672gat);
assign n971gat = ~(n111gat | n2840gat);
assign n247gat = ~(n334gat | n387gat | n330gat);
assign n145gat = ~(n144gat | n325gat);
assign n143gat = ~(n326gat | n247gat);
assign n970gat = ~(n372gat | n878gat);
assign n968gat = ~(n2789gat | n219gat);
assign n772gat = ~(n111gat | n2842gat);
assign n142gat = ~(n382gat | n326gat | n144gat);
assign n40gat = ~(n325gat | n383gat);
assign n39gat = ~(n383gat | n247gat);
assign n451gat = ~(n134gat | n372gat);
assign n446gat = ~(n219gat | n2781gat);
assign n139gat = ~(n253gat | n151gat | n254gat);
assign n136gat = ~(n253gat | n154gat);
assign n391gat = ~(n252gat | n468gat);
assign n390gat = ~(n469gat | n2877gat);
assign n1083gat = ~(n381gat | n375gat);
assign n1077gat = ~(n110gat | n2672gat);
assign n140gat = ~(n151gat | n253gat | n155gat);
assign n242gat = ~(n254gat | n241gat);
assign n240gat = ~(n255gat | n140gat);
assign n871gat = ~(n802gat | n375gat);
assign n797gat = ~(n110gat | n2734gat);
assign n324gat = ~(n255gat | n146gat | n241gat);
assign n238gat = ~(n147gat | n254gat);
assign n237gat = ~(n140gat | n147gat);
assign n1082gat = ~(n375gat | n380gat);
assign n796gat = ~(n2731gat | n110gat);
assign n85gat = ~(n17gat | n294gat | n637gat);
assign n180gat = ~(n286gat | n188gat | n287gat);
assign n68gat = ~(n85gat | n180gat);
assign n186gat = ~(n189gat | n287gat | n288gat);
assign n357gat = ~(n2726gat | n2860gat);
assign n82gat = ~(n16gat | n295gat | n637gat);
assign n12gat = ~(n186gat | n82gat);
assign n1599gat = ~(n1691gat | n336gat);
assign n1613gat = ~(n1544gat | n1698gat);
assign n1756gat = ~(n2512gat | n1769gat | n1773gat);
assign n1586gat = ~(n1869gat | n1683gat);
assign n1755gat = ~(n1769gat | n1773gat | n2512gat);
assign n2538gat = ~(n2620gat | n2625gat | n2488gat);
assign n2483gat = ~(n2537gat | n2482gat | n2486gat);
assign n1391gat = ~(n1513gat | n2442gat);
assign n1471gat = ~(n1334gat | n1858gat | n1604gat);
assign n1469gat = ~(n1858gat | n1608gat);
assign n1472gat = ~(n1476gat | n1471gat | n1469gat);
assign n1927gat = ~(n1790gat | n1635gat);
assign n1470gat = ~(n1472gat | n1747gat);
assign n1402gat = ~(n1858gat | n1393gat | n1604gat);
assign n1400gat = ~(n1674gat | n1403gat);
assign n1567gat = ~(n1634gat | n1735gat);
assign n1399gat = ~(n1806gat | n1338gat | n1584gat);
assign n1564gat = ~(n1584gat | n1719gat | n1790gat | n1576gat);
assign n1600gat = ~(n1685gat | n1427gat);
assign n1519gat = ~(n1584gat | n1339gat | n1600gat);
assign n1397gat = ~(n1519gat | n1401gat);
assign n1398gat = ~(n1455gat | n1397gat);
assign n2008gat = ~(n2012gat | n1774gat);
assign n2005gat = ~(n2002gat | n2857gat);
assign n1818gat = ~(n1823gat | n2005gat);
assign n1759gat = ~(n1818gat | n1935gat | n2765gat);
assign n1686gat = ~(n1774gat | n1869gat | n1684gat);
assign n1533gat = ~(n1524gat | n1403gat);
assign n1863gat = ~(n1991gat | n2283gat | n1989gat);
assign n1860gat = ~(n1988gat | n2216gat | n1862gat);
assign n1915gat = ~(n1859gat | n1919gat);
assign n1510gat = ~(n1584gat | n1460gat);
assign n1800gat = ~(n1635gat | n1919gat);
assign n1459gat = ~(n1595gat | n1454gat);
assign n1458gat = ~(n1510gat | n1459gat);
assign n1532gat = ~(n1677gat | n1458gat);
assign n1467gat = ~(n2289gat | n1468gat);
assign n1466gat = ~(n1392gat | n1461gat | n1396gat);
assign n1531gat = ~(n1507gat | n1477gat);
assign n1593gat = ~(n1551gat | n1310gat);
assign n1602gat = ~(n1594gat | n1587gat | n2989gat);
assign n1761gat = ~(n2985gat | n1602gat | n1681gat);
assign n1760gat = ~(n1681gat | n1602gat | n2985gat);
assign n1721gat = ~(n2442gat | n1690gat | n1978gat);
assign n520gat = ~(n374gat | n2862gat);
assign n519gat = ~(n2854gat | n374gat);
assign n518gat = ~(n520gat | n519gat);
assign n418gat = ~(n374gat | n2723gat);
assign n411gat = ~(n374gat | n2726gat);
assign n522gat = ~(n374gat | n2859gat);
assign n516gat = ~(n374gat | n2715gat);
assign n410gat = ~(n417gat | n413gat | n412gat | n406gat);
assign n354gat = ~(n411gat | n522gat);
assign n355gat = ~(n517gat | n410gat | n354gat);
assign n408gat = ~(n516gat | n407gat);
assign n526gat = ~(n2859gat | n740gat);
assign n531gat = ~(n740gat | n2854gat);
assign n530gat = ~(n2862gat | n740gat);
assign n525gat = ~(n526gat | n531gat | n530gat);
assign n356gat = ~(n2726gat | n740gat);
assign n415gat = ~(n2723gat | n740gat);
assign n521gat = ~(n740gat | n2715gat);
assign n532gat = ~(n527gat | n416gat | n528gat);
assign n359gat = ~(n290gat | n358gat);
assign n420gat = ~(n408gat | n359gat);
assign n523gat = ~(n522gat | n356gat);
assign n634gat = ~(n418gat | n521gat);
assign n414gat = ~(n411gat | n415gat);
assign n635gat = ~(n639gat | n634gat | n414gat);
assign n1100gat = ~(n1297gat | n1111gat);
assign n630gat = ~(n634gat | n523gat | n524gat);
assign n994gat = ~(n1112gat | n882gat);
assign n629gat = ~(n414gat | n634gat | n523gat);
assign n989gat = ~(n721gat | n741gat);
assign n632gat = ~(n414gat | n523gat | n633gat);
assign n880gat = ~(n926gat | n566gat);
assign n636gat = ~(n414gat | n633gat | n639gat);
assign n801gat = ~(n672gat | n670gat);
assign n879gat = ~(n2931gat | n801gat);
assign n1003gat = ~(n420gat | n879gat);
assign n1255gat = ~(n1123gat | n1225gat);
assign n1012gat = ~(n1007gat | n918gat);
assign n905gat = ~(n625gat | n1006gat);
assign n1009gat = ~(n1255gat | n2943gat);
assign n409gat = ~(n406gat | n407gat);
assign n292gat = ~(n415gat | n356gat);
assign n291gat = ~(n290gat | n292gat);
assign n419gat = ~(n409gat | n291gat);
assign n902gat = ~(n1009gat | n419gat);
assign n1099gat = ~(n1111gat | n1293gat);
assign n998gat = ~(n725gat | n741gat);
assign n995gat = ~(n823gat | n1112gat);
assign n980gat = ~(n875gat | n926gat);
assign n1001gat = ~(n420gat | n1002gat);
assign n1175gat = ~(n621gat | n1006gat);
assign n1174gat = ~(n845gat | n1007gat);
assign n1243gat = ~(n1281gat | n1123gat);
assign n1171gat = ~(n2960gat | n1243gat);
assign n999gat = ~(n419gat | n1171gat);
assign n1244gat = ~(n1123gat | n1134gat);
assign n1323gat = ~(n1007gat | n401gat);
assign n1264gat = ~(n1006gat | n617gat);
assign n1265gat = ~(n1244gat | n2969gat);
assign n892gat = ~(n419gat | n1265gat);
assign n981gat = ~(n926gat | n873gat);
assign n890gat = ~(n741gat | n702gat);
assign n889gat = ~(n1111gat | n1079gat);
assign n886gat = ~(n683gat | n1112gat);
assign n891gat = ~(n420gat | n888gat);
assign n904gat = ~(n1006gat | n490gat);
assign n903gat = ~(n1007gat | n397gat);
assign n1254gat = ~(n1123gat | n1044gat);
assign n1008gat = ~(n2942gat | n1254gat);
assign n900gat = ~(n419gat | n1008gat);
assign n1152gat = ~(n926gat | n1150gat);
assign n1092gat = ~(n1147gat | n1111gat);
assign n997gat = ~(n741gat | n393gat);
assign n993gat = ~(n1112gat | n698gat);
assign n895gat = ~(n420gat | n898gat);
assign n1094gat = ~(n1112gat | n583gat);
assign n1093gat = ~(n1111gat | n864gat);
assign n988gat = ~(n340gat | n741gat);
assign n984gat = ~(n926gat | n983gat);
assign n1178gat = ~(n420gat | n1179gat);
assign n1267gat = ~(n613gat | n1006gat);
assign n1257gat = ~(n1007gat | n274gat);
assign n1253gat = ~(n930gat | n1123gat);
assign n1266gat = ~(n2965gat | n1253gat);
assign n1116gat = ~(n419gat | n1266gat);
assign n1375gat = ~(n1006gat | n706gat);
assign n1324gat = ~(n164gat | n1007gat);
assign n1200gat = ~(n1120gat | n1123gat);
assign n1172gat = ~(n2961gat | n1200gat);
assign n899gat = ~(n419gat | n1172gat);
assign n1091gat = ~(n1111gat | n956gat);
assign n1088gat = ~(n1085gat | n926gat);
assign n992gat = ~(n815gat | n1112gat);
assign n987gat = ~(n741gat | n159gat);
assign n896gat = ~(n897gat | n420gat);
assign n1262gat = ~(n837gat | n1006gat);
assign n1260gat = ~(n1007gat | n278gat);
assign n1251gat = ~(n1123gat | n1071gat);
assign n1259gat = ~(n2967gat | n1251gat);
assign n901gat = ~(n419gat | n1259gat);
assign n1098gat = ~(n336gat | n741gat);
assign n1090gat = ~(n1111gat | n860gat);
assign n986gat = ~(n985gat | n926gat);
assign n885gat = ~(n579gat | n1112gat);
assign n893gat = ~(n894gat | n420gat);
assign n1097gat = ~(n270gat | n741gat);
assign n1089gat = ~(n1067gat | n1111gat);
assign n1087gat = ~(n926gat | n1084gat);
assign n991gat = ~(n1112gat | n679gat);
assign n1177gat = ~(n1180gat | n420gat);
assign n1212gat = ~(n1123gat | n1034gat);
assign n1326gat = ~(n1007gat | n282gat);
assign n1261gat = ~(n833gat | n1006gat);
assign n1263gat = ~(n1212gat | n2968gat);
assign n1115gat = ~(n1263gat | n419gat);
assign n977gat = ~(n670gat | n671gat);
assign n631gat = ~(n523gat | n633gat | n524gat);
assign n1096gat = ~(n819gat | n1112gat);
assign n1095gat = ~(n1240gat | n1111gat);
assign n990gat = ~(n841gat | n741gat);
assign n979gat = ~(n1601gat | n926gat);
assign n978gat = ~(n2944gat | n2945gat);
assign n1004gat = ~(n978gat | n420gat);
assign n1199gat = ~(n1123gat | n1284gat);
assign n1176gat = ~(n829gat | n1006gat);
assign n1173gat = ~(n1007gat | n1025gat);
assign n1252gat = ~(n1199gat | n2962gat);
assign n1000gat = ~(n419gat | n1252gat);
assign n1029gat = ~(n978gat | n455gat);
assign n1028gat = ~(n455gat | n879gat);
assign n1031gat = ~(n1002gat | n455gat);
assign n1030gat = ~(n455gat | n888gat);
assign n1011gat = ~(n455gat | n898gat);
assign n1181gat = ~(n455gat | n1179gat);
assign n1010gat = ~(n897gat | n455gat);
assign n1005gat = ~(n894gat | n455gat);
assign n1182gat = ~(n1180gat | n455gat);
assign n1757gat = ~(n1773gat | n1769gat);
assign n1745gat = ~(n1869gat | n1757gat);
assign n73gat = ~(n67gat | n2784gat);
assign n70gat = ~(n71gat | n2720gat);
assign n77gat = ~(n76gat | n2784gat);
assign n13gat = ~(n2720gat | n14gat);

endmodule
